module collision1
	(
		x,
		y,
		out
	);
	input 	[6:0]	x;
	input	[6:0] 	y;
	output 	[1:0]	out;
	wire [14:0] location;
	
	wire [19200: 0] COL;
assign COL[1] = 1'b1;
assign COL[2] = 1'b1;
assign COL[3] = 1'b1;
assign COL[4] = 1'b1;
assign COL[5] = 1'b1;
assign COL[6] = 1'b1;
assign COL[7] = 1'b1;
assign COL[8] = 1'b1;
assign COL[9] = 1'b1;
assign COL[10] = 1'b1;
assign COL[11] = 1'b1;
assign COL[12] = 1'b1;
assign COL[13] = 1'b1;
assign COL[14] = 1'b1;
assign COL[15] = 1'b1;
assign COL[16] = 1'b1;
assign COL[17] = 1'b1;
assign COL[18] = 1'b1;
assign COL[19] = 1'b1;
assign COL[20] = 1'b1;
assign COL[21] = 1'b1;
assign COL[22] = 1'b1;
assign COL[23] = 1'b1;
assign COL[24] = 1'b1;
assign COL[25] = 1'b1;
assign COL[26] = 1'b1;
assign COL[27] = 1'b1;
assign COL[28] = 1'b1;
assign COL[29] = 1'b1;
assign COL[30] = 1'b1;
assign COL[31] = 1'b1;
assign COL[32] = 1'b1;
assign COL[33] = 1'b1;
assign COL[34] = 1'b1;
assign COL[35] = 1'b1;
assign COL[36] = 1'b1;
assign COL[37] = 1'b1;
assign COL[38] = 1'b1;
assign COL[39] = 1'b1;
assign COL[40] = 1'b1;
assign COL[41] = 1'b1;
assign COL[42] = 1'b1;
assign COL[43] = 1'b1;
assign COL[44] = 1'b1;
assign COL[45] = 1'b1;
assign COL[46] = 1'b1;
assign COL[47] = 1'b1;
assign COL[48] = 1'b1;
assign COL[49] = 1'b1;
assign COL[50] = 1'b1;
assign COL[51] = 1'b1;
assign COL[52] = 1'b1;
assign COL[53] = 1'b1;
assign COL[54] = 1'b1;
assign COL[55] = 1'b1;
assign COL[56] = 1'b1;
assign COL[57] = 1'b1;
assign COL[58] = 1'b1;
assign COL[59] = 1'b1;
assign COL[60] = 1'b1;
assign COL[61] = 1'b1;
assign COL[62] = 1'b1;
assign COL[63] = 1'b1;
assign COL[64] = 1'b1;
assign COL[65] = 1'b1;
assign COL[66] = 1'b1;
assign COL[67] = 1'b1;
assign COL[68] = 1'b1;
assign COL[69] = 1'b1;
assign COL[70] = 1'b1;
assign COL[71] = 1'b1;
assign COL[72] = 1'b1;
assign COL[73] = 1'b1;
assign COL[74] = 1'b1;
assign COL[75] = 1'b1;
assign COL[76] = 1'b1;
assign COL[77] = 1'b1;
assign COL[78] = 1'b1;
assign COL[79] = 1'b1;
assign COL[80] = 1'b1;
assign COL[81] = 1'b1;
assign COL[82] = 1'b1;
assign COL[83] = 1'b1;
assign COL[84] = 1'b1;
assign COL[85] = 1'b1;
assign COL[86] = 1'b1;
assign COL[87] = 1'b1;
assign COL[88] = 1'b1;
assign COL[89] = 1'b1;
assign COL[90] = 1'b1;
assign COL[91] = 1'b1;
assign COL[92] = 1'b1;
assign COL[93] = 1'b1;
assign COL[94] = 1'b1;
assign COL[95] = 1'b0;
assign COL[96] = 1'b0;
assign COL[97] = 1'b0;
assign COL[98] = 1'b0;
assign COL[99] = 1'b0;
assign COL[100] = 1'b0;
assign COL[101] = 1'b0;
assign COL[102] = 1'b0;
assign COL[103] = 1'b0;
assign COL[104] = 1'b0;
assign COL[105] = 1'b0;
assign COL[106] = 1'b0;
assign COL[107] = 1'b0;
assign COL[108] = 1'b0;
assign COL[109] = 1'b0;
assign COL[110] = 1'b0;
assign COL[111] = 1'b0;
assign COL[112] = 1'b0;
assign COL[113] = 1'b0;
assign COL[114] = 1'b0;
assign COL[115] = 1'b0;
assign COL[116] = 1'b0;
assign COL[117] = 1'b0;
assign COL[118] = 1'b0;
assign COL[119] = 1'b0;
assign COL[120] = 1'b0;
assign COL[121] = 1'b0;
assign COL[122] = 1'b0;
assign COL[123] = 1'b0;
assign COL[124] = 1'b0;
assign COL[125] = 1'b0;
assign COL[126] = 1'b0;
assign COL[127] = 1'b0;
assign COL[128] = 1'b0;
assign COL[129] = 1'b0;
assign COL[130] = 1'b0;
assign COL[131] = 1'b0;
assign COL[132] = 1'b0;
assign COL[133] = 1'b0;
assign COL[134] = 1'b0;
assign COL[135] = 1'b0;
assign COL[136] = 1'b0;
assign COL[137] = 1'b0;
assign COL[138] = 1'b0;
assign COL[139] = 1'b0;
assign COL[140] = 1'b0;
assign COL[141] = 1'b0;
assign COL[142] = 1'b0;
assign COL[143] = 1'b0;
assign COL[144] = 1'b0;
assign COL[145] = 1'b0;
assign COL[146] = 1'b0;
assign COL[147] = 1'b0;
assign COL[148] = 1'b0;
assign COL[149] = 1'b0;
assign COL[150] = 1'b0;
assign COL[151] = 1'b0;
assign COL[152] = 1'b0;
assign COL[153] = 1'b0;
assign COL[154] = 1'b0;
assign COL[155] = 1'b0;
assign COL[156] = 1'b0;
assign COL[157] = 1'b0;
assign COL[158] = 1'b0;
assign COL[159] = 1'b0;
assign COL[160] = 1'b0;
assign COL[161] = 1'b1;
assign COL[162] = 1'b1;
assign COL[163] = 1'b1;
assign COL[164] = 1'b1;
assign COL[165] = 1'b1;
assign COL[166] = 1'b1;
assign COL[167] = 1'b1;
assign COL[168] = 1'b1;
assign COL[169] = 1'b1;
assign COL[170] = 1'b1;
assign COL[171] = 1'b1;
assign COL[172] = 1'b1;
assign COL[173] = 1'b1;
assign COL[174] = 1'b1;
assign COL[175] = 1'b1;
assign COL[176] = 1'b1;
assign COL[177] = 1'b1;
assign COL[178] = 1'b1;
assign COL[179] = 1'b1;
assign COL[180] = 1'b1;
assign COL[181] = 1'b1;
assign COL[182] = 1'b1;
assign COL[183] = 1'b1;
assign COL[184] = 1'b1;
assign COL[185] = 1'b1;
assign COL[186] = 1'b1;
assign COL[187] = 1'b1;
assign COL[188] = 1'b1;
assign COL[189] = 1'b1;
assign COL[190] = 1'b1;
assign COL[191] = 1'b1;
assign COL[192] = 1'b1;
assign COL[193] = 1'b1;
assign COL[194] = 1'b1;
assign COL[195] = 1'b1;
assign COL[196] = 1'b1;
assign COL[197] = 1'b1;
assign COL[198] = 1'b1;
assign COL[199] = 1'b1;
assign COL[200] = 1'b1;
assign COL[201] = 1'b1;
assign COL[202] = 1'b1;
assign COL[203] = 1'b1;
assign COL[204] = 1'b1;
assign COL[205] = 1'b1;
assign COL[206] = 1'b1;
assign COL[207] = 1'b1;
assign COL[208] = 1'b1;
assign COL[209] = 1'b1;
assign COL[210] = 1'b1;
assign COL[211] = 1'b1;
assign COL[212] = 1'b1;
assign COL[213] = 1'b1;
assign COL[214] = 1'b1;
assign COL[215] = 1'b1;
assign COL[216] = 1'b1;
assign COL[217] = 1'b1;
assign COL[218] = 1'b1;
assign COL[219] = 1'b1;
assign COL[220] = 1'b1;
assign COL[221] = 1'b1;
assign COL[222] = 1'b1;
assign COL[223] = 1'b1;
assign COL[224] = 1'b1;
assign COL[225] = 1'b1;
assign COL[226] = 1'b1;
assign COL[227] = 1'b1;
assign COL[228] = 1'b1;
assign COL[229] = 1'b1;
assign COL[230] = 1'b1;
assign COL[231] = 1'b1;
assign COL[232] = 1'b1;
assign COL[233] = 1'b1;
assign COL[234] = 1'b1;
assign COL[235] = 1'b1;
assign COL[236] = 1'b1;
assign COL[237] = 1'b1;
assign COL[238] = 1'b1;
assign COL[239] = 1'b1;
assign COL[240] = 1'b1;
assign COL[241] = 1'b1;
assign COL[242] = 1'b1;
assign COL[243] = 1'b1;
assign COL[244] = 1'b1;
assign COL[245] = 1'b1;
assign COL[246] = 1'b1;
assign COL[247] = 1'b1;
assign COL[248] = 1'b1;
assign COL[249] = 1'b1;
assign COL[250] = 1'b1;
assign COL[251] = 1'b1;
assign COL[252] = 1'b1;
assign COL[253] = 1'b1;
assign COL[254] = 1'b1;
assign COL[255] = 1'b0;
assign COL[256] = 1'b0;
assign COL[257] = 1'b0;
assign COL[258] = 1'b0;
assign COL[259] = 1'b0;
assign COL[260] = 1'b0;
assign COL[261] = 1'b0;
assign COL[262] = 1'b0;
assign COL[263] = 1'b0;
assign COL[264] = 1'b0;
assign COL[265] = 1'b0;
assign COL[266] = 1'b0;
assign COL[267] = 1'b0;
assign COL[268] = 1'b0;
assign COL[269] = 1'b0;
assign COL[270] = 1'b0;
assign COL[271] = 1'b0;
assign COL[272] = 1'b0;
assign COL[273] = 1'b0;
assign COL[274] = 1'b0;
assign COL[275] = 1'b0;
assign COL[276] = 1'b0;
assign COL[277] = 1'b0;
assign COL[278] = 1'b0;
assign COL[279] = 1'b0;
assign COL[280] = 1'b0;
assign COL[281] = 1'b0;
assign COL[282] = 1'b0;
assign COL[283] = 1'b0;
assign COL[284] = 1'b0;
assign COL[285] = 1'b0;
assign COL[286] = 1'b0;
assign COL[287] = 1'b0;
assign COL[288] = 1'b0;
assign COL[289] = 1'b0;
assign COL[290] = 1'b0;
assign COL[291] = 1'b0;
assign COL[292] = 1'b0;
assign COL[293] = 1'b0;
assign COL[294] = 1'b0;
assign COL[295] = 1'b0;
assign COL[296] = 1'b0;
assign COL[297] = 1'b0;
assign COL[298] = 1'b0;
assign COL[299] = 1'b0;
assign COL[300] = 1'b0;
assign COL[301] = 1'b0;
assign COL[302] = 1'b0;
assign COL[303] = 1'b0;
assign COL[304] = 1'b0;
assign COL[305] = 1'b0;
assign COL[306] = 1'b0;
assign COL[307] = 1'b0;
assign COL[308] = 1'b0;
assign COL[309] = 1'b0;
assign COL[310] = 1'b0;
assign COL[311] = 1'b0;
assign COL[312] = 1'b0;
assign COL[313] = 1'b0;
assign COL[314] = 1'b0;
assign COL[315] = 1'b0;
assign COL[316] = 1'b0;
assign COL[317] = 1'b0;
assign COL[318] = 1'b0;
assign COL[319] = 1'b0;
assign COL[320] = 1'b0;
assign COL[321] = 1'b1;
assign COL[322] = 1'b1;
assign COL[323] = 1'b1;
assign COL[324] = 1'b1;
assign COL[325] = 1'b1;
assign COL[326] = 1'b1;
assign COL[327] = 1'b1;
assign COL[328] = 1'b1;
assign COL[329] = 1'b1;
assign COL[330] = 1'b1;
assign COL[331] = 1'b1;
assign COL[332] = 1'b1;
assign COL[333] = 1'b1;
assign COL[334] = 1'b1;
assign COL[335] = 1'b1;
assign COL[336] = 1'b1;
assign COL[337] = 1'b1;
assign COL[338] = 1'b1;
assign COL[339] = 1'b1;
assign COL[340] = 1'b1;
assign COL[341] = 1'b1;
assign COL[342] = 1'b1;
assign COL[343] = 1'b1;
assign COL[344] = 1'b1;
assign COL[345] = 1'b1;
assign COL[346] = 1'b1;
assign COL[347] = 1'b1;
assign COL[348] = 1'b1;
assign COL[349] = 1'b1;
assign COL[350] = 1'b1;
assign COL[351] = 1'b1;
assign COL[352] = 1'b1;
assign COL[353] = 1'b1;
assign COL[354] = 1'b1;
assign COL[355] = 1'b1;
assign COL[356] = 1'b1;
assign COL[357] = 1'b1;
assign COL[358] = 1'b1;
assign COL[359] = 1'b1;
assign COL[360] = 1'b1;
assign COL[361] = 1'b1;
assign COL[362] = 1'b1;
assign COL[363] = 1'b1;
assign COL[364] = 1'b1;
assign COL[365] = 1'b1;
assign COL[366] = 1'b1;
assign COL[367] = 1'b1;
assign COL[368] = 1'b1;
assign COL[369] = 1'b1;
assign COL[370] = 1'b1;
assign COL[371] = 1'b1;
assign COL[372] = 1'b1;
assign COL[373] = 1'b1;
assign COL[374] = 1'b1;
assign COL[375] = 1'b1;
assign COL[376] = 1'b1;
assign COL[377] = 1'b1;
assign COL[378] = 1'b1;
assign COL[379] = 1'b1;
assign COL[380] = 1'b1;
assign COL[381] = 1'b1;
assign COL[382] = 1'b1;
assign COL[383] = 1'b1;
assign COL[384] = 1'b1;
assign COL[385] = 1'b1;
assign COL[386] = 1'b1;
assign COL[387] = 1'b1;
assign COL[388] = 1'b1;
assign COL[389] = 1'b1;
assign COL[390] = 1'b1;
assign COL[391] = 1'b1;
assign COL[392] = 1'b1;
assign COL[393] = 1'b1;
assign COL[394] = 1'b1;
assign COL[395] = 1'b1;
assign COL[396] = 1'b1;
assign COL[397] = 1'b1;
assign COL[398] = 1'b1;
assign COL[399] = 1'b1;
assign COL[400] = 1'b1;
assign COL[401] = 1'b1;
assign COL[402] = 1'b1;
assign COL[403] = 1'b1;
assign COL[404] = 1'b1;
assign COL[405] = 1'b1;
assign COL[406] = 1'b1;
assign COL[407] = 1'b1;
assign COL[408] = 1'b1;
assign COL[409] = 1'b1;
assign COL[410] = 1'b1;
assign COL[411] = 1'b1;
assign COL[412] = 1'b1;
assign COL[413] = 1'b1;
assign COL[414] = 1'b1;
assign COL[415] = 1'b0;
assign COL[416] = 1'b0;
assign COL[417] = 1'b0;
assign COL[418] = 1'b0;
assign COL[419] = 1'b0;
assign COL[420] = 1'b0;
assign COL[421] = 1'b0;
assign COL[422] = 1'b0;
assign COL[423] = 1'b0;
assign COL[424] = 1'b0;
assign COL[425] = 1'b0;
assign COL[426] = 1'b0;
assign COL[427] = 1'b0;
assign COL[428] = 1'b0;
assign COL[429] = 1'b0;
assign COL[430] = 1'b0;
assign COL[431] = 1'b0;
assign COL[432] = 1'b0;
assign COL[433] = 1'b0;
assign COL[434] = 1'b0;
assign COL[435] = 1'b0;
assign COL[436] = 1'b0;
assign COL[437] = 1'b0;
assign COL[438] = 1'b0;
assign COL[439] = 1'b0;
assign COL[440] = 1'b0;
assign COL[441] = 1'b0;
assign COL[442] = 1'b0;
assign COL[443] = 1'b0;
assign COL[444] = 1'b0;
assign COL[445] = 1'b0;
assign COL[446] = 1'b0;
assign COL[447] = 1'b0;
assign COL[448] = 1'b0;
assign COL[449] = 1'b0;
assign COL[450] = 1'b0;
assign COL[451] = 1'b0;
assign COL[452] = 1'b0;
assign COL[453] = 1'b0;
assign COL[454] = 1'b0;
assign COL[455] = 1'b0;
assign COL[456] = 1'b0;
assign COL[457] = 1'b0;
assign COL[458] = 1'b0;
assign COL[459] = 1'b0;
assign COL[460] = 1'b0;
assign COL[461] = 1'b0;
assign COL[462] = 1'b0;
assign COL[463] = 1'b0;
assign COL[464] = 1'b0;
assign COL[465] = 1'b0;
assign COL[466] = 1'b0;
assign COL[467] = 1'b0;
assign COL[468] = 1'b0;
assign COL[469] = 1'b0;
assign COL[470] = 1'b0;
assign COL[471] = 1'b0;
assign COL[472] = 1'b0;
assign COL[473] = 1'b0;
assign COL[474] = 1'b0;
assign COL[475] = 1'b0;
assign COL[476] = 1'b0;
assign COL[477] = 1'b0;
assign COL[478] = 1'b0;
assign COL[479] = 1'b0;
assign COL[480] = 1'b0;
assign COL[481] = 1'b1;
assign COL[482] = 1'b1;
assign COL[483] = 1'b1;
assign COL[484] = 1'b1;
assign COL[485] = 1'b1;
assign COL[486] = 1'b1;
assign COL[487] = 1'b1;
assign COL[488] = 1'b1;
assign COL[489] = 1'b1;
assign COL[490] = 1'b1;
assign COL[491] = 1'b1;
assign COL[492] = 1'b1;
assign COL[493] = 1'b1;
assign COL[494] = 1'b1;
assign COL[495] = 1'b1;
assign COL[496] = 1'b1;
assign COL[497] = 1'b1;
assign COL[498] = 1'b1;
assign COL[499] = 1'b1;
assign COL[500] = 1'b1;
assign COL[501] = 1'b1;
assign COL[502] = 1'b1;
assign COL[503] = 1'b1;
assign COL[504] = 1'b1;
assign COL[505] = 1'b1;
assign COL[506] = 1'b1;
assign COL[507] = 1'b1;
assign COL[508] = 1'b1;
assign COL[509] = 1'b1;
assign COL[510] = 1'b1;
assign COL[511] = 1'b1;
assign COL[512] = 1'b1;
assign COL[513] = 1'b1;
assign COL[514] = 1'b1;
assign COL[515] = 1'b1;
assign COL[516] = 1'b1;
assign COL[517] = 1'b1;
assign COL[518] = 1'b1;
assign COL[519] = 1'b1;
assign COL[520] = 1'b1;
assign COL[521] = 1'b1;
assign COL[522] = 1'b1;
assign COL[523] = 1'b1;
assign COL[524] = 1'b1;
assign COL[525] = 1'b1;
assign COL[526] = 1'b1;
assign COL[527] = 1'b1;
assign COL[528] = 1'b1;
assign COL[529] = 1'b1;
assign COL[530] = 1'b1;
assign COL[531] = 1'b1;
assign COL[532] = 1'b1;
assign COL[533] = 1'b1;
assign COL[534] = 1'b1;
assign COL[535] = 1'b1;
assign COL[536] = 1'b1;
assign COL[537] = 1'b1;
assign COL[538] = 1'b1;
assign COL[539] = 1'b1;
assign COL[540] = 1'b1;
assign COL[541] = 1'b1;
assign COL[542] = 1'b1;
assign COL[543] = 1'b1;
assign COL[544] = 1'b1;
assign COL[545] = 1'b1;
assign COL[546] = 1'b1;
assign COL[547] = 1'b1;
assign COL[548] = 1'b1;
assign COL[549] = 1'b1;
assign COL[550] = 1'b1;
assign COL[551] = 1'b1;
assign COL[552] = 1'b1;
assign COL[553] = 1'b1;
assign COL[554] = 1'b1;
assign COL[555] = 1'b1;
assign COL[556] = 1'b1;
assign COL[557] = 1'b1;
assign COL[558] = 1'b1;
assign COL[559] = 1'b1;
assign COL[560] = 1'b1;
assign COL[561] = 1'b1;
assign COL[562] = 1'b1;
assign COL[563] = 1'b1;
assign COL[564] = 1'b1;
assign COL[565] = 1'b1;
assign COL[566] = 1'b1;
assign COL[567] = 1'b1;
assign COL[568] = 1'b1;
assign COL[569] = 1'b1;
assign COL[570] = 1'b1;
assign COL[571] = 1'b1;
assign COL[572] = 1'b1;
assign COL[573] = 1'b1;
assign COL[574] = 1'b1;
assign COL[575] = 1'b0;
assign COL[576] = 1'b0;
assign COL[577] = 1'b0;
assign COL[578] = 1'b0;
assign COL[579] = 1'b0;
assign COL[580] = 1'b0;
assign COL[581] = 1'b0;
assign COL[582] = 1'b0;
assign COL[583] = 1'b0;
assign COL[584] = 1'b0;
assign COL[585] = 1'b0;
assign COL[586] = 1'b0;
assign COL[587] = 1'b0;
assign COL[588] = 1'b0;
assign COL[589] = 1'b0;
assign COL[590] = 1'b0;
assign COL[591] = 1'b0;
assign COL[592] = 1'b0;
assign COL[593] = 1'b0;
assign COL[594] = 1'b0;
assign COL[595] = 1'b0;
assign COL[596] = 1'b0;
assign COL[597] = 1'b0;
assign COL[598] = 1'b0;
assign COL[599] = 1'b0;
assign COL[600] = 1'b0;
assign COL[601] = 1'b0;
assign COL[602] = 1'b0;
assign COL[603] = 1'b0;
assign COL[604] = 1'b0;
assign COL[605] = 1'b0;
assign COL[606] = 1'b0;
assign COL[607] = 1'b0;
assign COL[608] = 1'b0;
assign COL[609] = 1'b0;
assign COL[610] = 1'b0;
assign COL[611] = 1'b0;
assign COL[612] = 1'b0;
assign COL[613] = 1'b0;
assign COL[614] = 1'b0;
assign COL[615] = 1'b0;
assign COL[616] = 1'b0;
assign COL[617] = 1'b0;
assign COL[618] = 1'b0;
assign COL[619] = 1'b0;
assign COL[620] = 1'b0;
assign COL[621] = 1'b0;
assign COL[622] = 1'b0;
assign COL[623] = 1'b0;
assign COL[624] = 1'b0;
assign COL[625] = 1'b0;
assign COL[626] = 1'b0;
assign COL[627] = 1'b0;
assign COL[628] = 1'b0;
assign COL[629] = 1'b0;
assign COL[630] = 1'b0;
assign COL[631] = 1'b0;
assign COL[632] = 1'b0;
assign COL[633] = 1'b0;
assign COL[634] = 1'b0;
assign COL[635] = 1'b0;
assign COL[636] = 1'b0;
assign COL[637] = 1'b0;
assign COL[638] = 1'b0;
assign COL[639] = 1'b0;
assign COL[640] = 1'b0;
assign COL[641] = 1'b1;
assign COL[642] = 1'b1;
assign COL[643] = 1'b1;
assign COL[644] = 1'b1;
assign COL[645] = 1'b1;
assign COL[646] = 1'b1;
assign COL[647] = 1'b1;
assign COL[648] = 1'b1;
assign COL[649] = 1'b1;
assign COL[650] = 1'b1;
assign COL[651] = 1'b1;
assign COL[652] = 1'b1;
assign COL[653] = 1'b1;
assign COL[654] = 1'b1;
assign COL[655] = 1'b1;
assign COL[656] = 1'b1;
assign COL[657] = 1'b1;
assign COL[658] = 1'b1;
assign COL[659] = 1'b1;
assign COL[660] = 1'b1;
assign COL[661] = 1'b1;
assign COL[662] = 1'b1;
assign COL[663] = 1'b1;
assign COL[664] = 1'b1;
assign COL[665] = 1'b1;
assign COL[666] = 1'b1;
assign COL[667] = 1'b1;
assign COL[668] = 1'b1;
assign COL[669] = 1'b1;
assign COL[670] = 1'b1;
assign COL[671] = 1'b1;
assign COL[672] = 1'b1;
assign COL[673] = 1'b1;
assign COL[674] = 1'b1;
assign COL[675] = 1'b1;
assign COL[676] = 1'b1;
assign COL[677] = 1'b1;
assign COL[678] = 1'b1;
assign COL[679] = 1'b1;
assign COL[680] = 1'b1;
assign COL[681] = 1'b1;
assign COL[682] = 1'b1;
assign COL[683] = 1'b1;
assign COL[684] = 1'b1;
assign COL[685] = 1'b1;
assign COL[686] = 1'b1;
assign COL[687] = 1'b1;
assign COL[688] = 1'b1;
assign COL[689] = 1'b1;
assign COL[690] = 1'b1;
assign COL[691] = 1'b1;
assign COL[692] = 1'b1;
assign COL[693] = 1'b1;
assign COL[694] = 1'b1;
assign COL[695] = 1'b1;
assign COL[696] = 1'b1;
assign COL[697] = 1'b1;
assign COL[698] = 1'b1;
assign COL[699] = 1'b1;
assign COL[700] = 1'b1;
assign COL[701] = 1'b1;
assign COL[702] = 1'b1;
assign COL[703] = 1'b1;
assign COL[704] = 1'b1;
assign COL[705] = 1'b1;
assign COL[706] = 1'b1;
assign COL[707] = 1'b1;
assign COL[708] = 1'b1;
assign COL[709] = 1'b1;
assign COL[710] = 1'b1;
assign COL[711] = 1'b1;
assign COL[712] = 1'b1;
assign COL[713] = 1'b1;
assign COL[714] = 1'b1;
assign COL[715] = 1'b1;
assign COL[716] = 1'b1;
assign COL[717] = 1'b1;
assign COL[718] = 1'b1;
assign COL[719] = 1'b1;
assign COL[720] = 1'b1;
assign COL[721] = 1'b1;
assign COL[722] = 1'b1;
assign COL[723] = 1'b1;
assign COL[724] = 1'b1;
assign COL[725] = 1'b1;
assign COL[726] = 1'b1;
assign COL[727] = 1'b1;
assign COL[728] = 1'b1;
assign COL[729] = 1'b1;
assign COL[730] = 1'b1;
assign COL[731] = 1'b1;
assign COL[732] = 1'b1;
assign COL[733] = 1'b1;
assign COL[734] = 1'b1;
assign COL[735] = 1'b0;
assign COL[736] = 1'b0;
assign COL[737] = 1'b0;
assign COL[738] = 1'b0;
assign COL[739] = 1'b0;
assign COL[740] = 1'b0;
assign COL[741] = 1'b0;
assign COL[742] = 1'b0;
assign COL[743] = 1'b0;
assign COL[744] = 1'b0;
assign COL[745] = 1'b0;
assign COL[746] = 1'b0;
assign COL[747] = 1'b0;
assign COL[748] = 1'b0;
assign COL[749] = 1'b0;
assign COL[750] = 1'b0;
assign COL[751] = 1'b0;
assign COL[752] = 1'b0;
assign COL[753] = 1'b0;
assign COL[754] = 1'b0;
assign COL[755] = 1'b0;
assign COL[756] = 1'b0;
assign COL[757] = 1'b0;
assign COL[758] = 1'b0;
assign COL[759] = 1'b0;
assign COL[760] = 1'b0;
assign COL[761] = 1'b0;
assign COL[762] = 1'b0;
assign COL[763] = 1'b0;
assign COL[764] = 1'b0;
assign COL[765] = 1'b0;
assign COL[766] = 1'b0;
assign COL[767] = 1'b0;
assign COL[768] = 1'b0;
assign COL[769] = 1'b0;
assign COL[770] = 1'b0;
assign COL[771] = 1'b0;
assign COL[772] = 1'b0;
assign COL[773] = 1'b0;
assign COL[774] = 1'b0;
assign COL[775] = 1'b0;
assign COL[776] = 1'b0;
assign COL[777] = 1'b0;
assign COL[778] = 1'b0;
assign COL[779] = 1'b0;
assign COL[780] = 1'b0;
assign COL[781] = 1'b0;
assign COL[782] = 1'b0;
assign COL[783] = 1'b0;
assign COL[784] = 1'b0;
assign COL[785] = 1'b0;
assign COL[786] = 1'b0;
assign COL[787] = 1'b0;
assign COL[788] = 1'b0;
assign COL[789] = 1'b0;
assign COL[790] = 1'b0;
assign COL[791] = 1'b0;
assign COL[792] = 1'b0;
assign COL[793] = 1'b0;
assign COL[794] = 1'b0;
assign COL[795] = 1'b0;
assign COL[796] = 1'b0;
assign COL[797] = 1'b0;
assign COL[798] = 1'b0;
assign COL[799] = 1'b0;
assign COL[800] = 1'b0;
assign COL[801] = 1'b1;
assign COL[802] = 1'b1;
assign COL[803] = 1'b1;
assign COL[804] = 1'b1;
assign COL[805] = 1'b1;
assign COL[806] = 1'b0;
assign COL[807] = 1'b0;
assign COL[808] = 1'b0;
assign COL[809] = 1'b0;
assign COL[810] = 1'b0;
assign COL[811] = 1'b0;
assign COL[812] = 1'b0;
assign COL[813] = 1'b0;
assign COL[814] = 1'b0;
assign COL[815] = 1'b0;
assign COL[816] = 1'b0;
assign COL[817] = 1'b0;
assign COL[818] = 1'b0;
assign COL[819] = 1'b0;
assign COL[820] = 1'b0;
assign COL[821] = 1'b0;
assign COL[822] = 1'b0;
assign COL[823] = 1'b0;
assign COL[824] = 1'b0;
assign COL[825] = 1'b0;
assign COL[826] = 1'b0;
assign COL[827] = 1'b0;
assign COL[828] = 1'b0;
assign COL[829] = 1'b0;
assign COL[830] = 1'b0;
assign COL[831] = 1'b0;
assign COL[832] = 1'b0;
assign COL[833] = 1'b0;
assign COL[834] = 1'b0;
assign COL[835] = 1'b0;
assign COL[836] = 1'b0;
assign COL[837] = 1'b0;
assign COL[838] = 1'b0;
assign COL[839] = 1'b0;
assign COL[840] = 1'b1;
assign COL[841] = 1'b1;
assign COL[842] = 1'b1;
assign COL[843] = 1'b1;
assign COL[844] = 1'b0;
assign COL[845] = 1'b0;
assign COL[846] = 1'b0;
assign COL[847] = 1'b0;
assign COL[848] = 1'b0;
assign COL[849] = 1'b0;
assign COL[850] = 1'b0;
assign COL[851] = 1'b0;
assign COL[852] = 1'b0;
assign COL[853] = 1'b0;
assign COL[854] = 1'b0;
assign COL[855] = 1'b0;
assign COL[856] = 1'b0;
assign COL[857] = 1'b0;
assign COL[858] = 1'b0;
assign COL[859] = 1'b0;
assign COL[860] = 1'b0;
assign COL[861] = 1'b0;
assign COL[862] = 1'b0;
assign COL[863] = 1'b0;
assign COL[864] = 1'b0;
assign COL[865] = 1'b0;
assign COL[866] = 1'b0;
assign COL[867] = 1'b0;
assign COL[868] = 1'b0;
assign COL[869] = 1'b0;
assign COL[870] = 1'b0;
assign COL[871] = 1'b0;
assign COL[872] = 1'b1;
assign COL[873] = 1'b1;
assign COL[874] = 1'b1;
assign COL[875] = 1'b1;
assign COL[876] = 1'b0;
assign COL[877] = 1'b0;
assign COL[878] = 1'b0;
assign COL[879] = 1'b0;
assign COL[880] = 1'b0;
assign COL[881] = 1'b0;
assign COL[882] = 1'b0;
assign COL[883] = 1'b0;
assign COL[884] = 1'b0;
assign COL[885] = 1'b0;
assign COL[886] = 1'b0;
assign COL[887] = 1'b0;
assign COL[888] = 1'b0;
assign COL[889] = 1'b0;
assign COL[890] = 1'b1;
assign COL[891] = 1'b1;
assign COL[892] = 1'b1;
assign COL[893] = 1'b1;
assign COL[894] = 1'b1;
assign COL[895] = 1'b0;
assign COL[896] = 1'b0;
assign COL[897] = 1'b0;
assign COL[898] = 1'b0;
assign COL[899] = 1'b0;
assign COL[900] = 1'b0;
assign COL[901] = 1'b0;
assign COL[902] = 1'b0;
assign COL[903] = 1'b0;
assign COL[904] = 1'b0;
assign COL[905] = 1'b0;
assign COL[906] = 1'b0;
assign COL[907] = 1'b0;
assign COL[908] = 1'b0;
assign COL[909] = 1'b0;
assign COL[910] = 1'b0;
assign COL[911] = 1'b0;
assign COL[912] = 1'b0;
assign COL[913] = 1'b0;
assign COL[914] = 1'b0;
assign COL[915] = 1'b0;
assign COL[916] = 1'b0;
assign COL[917] = 1'b0;
assign COL[918] = 1'b0;
assign COL[919] = 1'b0;
assign COL[920] = 1'b0;
assign COL[921] = 1'b0;
assign COL[922] = 1'b0;
assign COL[923] = 1'b0;
assign COL[924] = 1'b0;
assign COL[925] = 1'b0;
assign COL[926] = 1'b0;
assign COL[927] = 1'b0;
assign COL[928] = 1'b0;
assign COL[929] = 1'b0;
assign COL[930] = 1'b0;
assign COL[931] = 1'b0;
assign COL[932] = 1'b0;
assign COL[933] = 1'b0;
assign COL[934] = 1'b0;
assign COL[935] = 1'b0;
assign COL[936] = 1'b0;
assign COL[937] = 1'b0;
assign COL[938] = 1'b0;
assign COL[939] = 1'b0;
assign COL[940] = 1'b0;
assign COL[941] = 1'b0;
assign COL[942] = 1'b0;
assign COL[943] = 1'b0;
assign COL[944] = 1'b0;
assign COL[945] = 1'b0;
assign COL[946] = 1'b0;
assign COL[947] = 1'b0;
assign COL[948] = 1'b0;
assign COL[949] = 1'b0;
assign COL[950] = 1'b0;
assign COL[951] = 1'b0;
assign COL[952] = 1'b0;
assign COL[953] = 1'b0;
assign COL[954] = 1'b0;
assign COL[955] = 1'b0;
assign COL[956] = 1'b0;
assign COL[957] = 1'b0;
assign COL[958] = 1'b0;
assign COL[959] = 1'b0;
assign COL[960] = 1'b0;
assign COL[961] = 1'b1;
assign COL[962] = 1'b1;
assign COL[963] = 1'b1;
assign COL[964] = 1'b1;
assign COL[965] = 1'b1;
assign COL[966] = 1'b0;
assign COL[967] = 1'b0;
assign COL[968] = 1'b0;
assign COL[969] = 1'b0;
assign COL[970] = 1'b0;
assign COL[971] = 1'b0;
assign COL[972] = 1'b0;
assign COL[973] = 1'b0;
assign COL[974] = 1'b0;
assign COL[975] = 1'b0;
assign COL[976] = 1'b0;
assign COL[977] = 1'b0;
assign COL[978] = 1'b0;
assign COL[979] = 1'b0;
assign COL[980] = 1'b0;
assign COL[981] = 1'b0;
assign COL[982] = 1'b0;
assign COL[983] = 1'b0;
assign COL[984] = 1'b0;
assign COL[985] = 1'b0;
assign COL[986] = 1'b0;
assign COL[987] = 1'b0;
assign COL[988] = 1'b0;
assign COL[989] = 1'b0;
assign COL[990] = 1'b0;
assign COL[991] = 1'b0;
assign COL[992] = 1'b0;
assign COL[993] = 1'b0;
assign COL[994] = 1'b0;
assign COL[995] = 1'b0;
assign COL[996] = 1'b0;
assign COL[997] = 1'b0;
assign COL[998] = 1'b0;
assign COL[999] = 1'b0;
assign COL[1000] = 1'b1;
assign COL[1001] = 1'b1;
assign COL[1002] = 1'b1;
assign COL[1003] = 1'b1;
assign COL[1004] = 1'b0;
assign COL[1005] = 1'b0;
assign COL[1006] = 1'b0;
assign COL[1007] = 1'b0;
assign COL[1008] = 1'b0;
assign COL[1009] = 1'b0;
assign COL[1010] = 1'b0;
assign COL[1011] = 1'b0;
assign COL[1012] = 1'b0;
assign COL[1013] = 1'b0;
assign COL[1014] = 1'b0;
assign COL[1015] = 1'b0;
assign COL[1016] = 1'b0;
assign COL[1017] = 1'b0;
assign COL[1018] = 1'b0;
assign COL[1019] = 1'b0;
assign COL[1020] = 1'b0;
assign COL[1021] = 1'b0;
assign COL[1022] = 1'b0;
assign COL[1023] = 1'b0;
assign COL[1024] = 1'b0;
assign COL[1025] = 1'b0;
assign COL[1026] = 1'b0;
assign COL[1027] = 1'b0;
assign COL[1028] = 1'b0;
assign COL[1029] = 1'b0;
assign COL[1030] = 1'b0;
assign COL[1031] = 1'b0;
assign COL[1032] = 1'b1;
assign COL[1033] = 1'b1;
assign COL[1034] = 1'b1;
assign COL[1035] = 1'b1;
assign COL[1036] = 1'b0;
assign COL[1037] = 1'b0;
assign COL[1038] = 1'b0;
assign COL[1039] = 1'b0;
assign COL[1040] = 1'b0;
assign COL[1041] = 1'b0;
assign COL[1042] = 1'b0;
assign COL[1043] = 1'b0;
assign COL[1044] = 1'b0;
assign COL[1045] = 1'b0;
assign COL[1046] = 1'b0;
assign COL[1047] = 1'b0;
assign COL[1048] = 1'b0;
assign COL[1049] = 1'b0;
assign COL[1050] = 1'b1;
assign COL[1051] = 1'b1;
assign COL[1052] = 1'b1;
assign COL[1053] = 1'b1;
assign COL[1054] = 1'b1;
assign COL[1055] = 1'b0;
assign COL[1056] = 1'b0;
assign COL[1057] = 1'b0;
assign COL[1058] = 1'b0;
assign COL[1059] = 1'b0;
assign COL[1060] = 1'b0;
assign COL[1061] = 1'b0;
assign COL[1062] = 1'b0;
assign COL[1063] = 1'b0;
assign COL[1064] = 1'b0;
assign COL[1065] = 1'b0;
assign COL[1066] = 1'b0;
assign COL[1067] = 1'b0;
assign COL[1068] = 1'b0;
assign COL[1069] = 1'b0;
assign COL[1070] = 1'b0;
assign COL[1071] = 1'b0;
assign COL[1072] = 1'b0;
assign COL[1073] = 1'b0;
assign COL[1074] = 1'b0;
assign COL[1075] = 1'b0;
assign COL[1076] = 1'b0;
assign COL[1077] = 1'b0;
assign COL[1078] = 1'b0;
assign COL[1079] = 1'b0;
assign COL[1080] = 1'b0;
assign COL[1081] = 1'b0;
assign COL[1082] = 1'b0;
assign COL[1083] = 1'b0;
assign COL[1084] = 1'b0;
assign COL[1085] = 1'b0;
assign COL[1086] = 1'b0;
assign COL[1087] = 1'b0;
assign COL[1088] = 1'b0;
assign COL[1089] = 1'b0;
assign COL[1090] = 1'b0;
assign COL[1091] = 1'b0;
assign COL[1092] = 1'b0;
assign COL[1093] = 1'b0;
assign COL[1094] = 1'b0;
assign COL[1095] = 1'b0;
assign COL[1096] = 1'b0;
assign COL[1097] = 1'b0;
assign COL[1098] = 1'b0;
assign COL[1099] = 1'b0;
assign COL[1100] = 1'b0;
assign COL[1101] = 1'b0;
assign COL[1102] = 1'b0;
assign COL[1103] = 1'b0;
assign COL[1104] = 1'b0;
assign COL[1105] = 1'b0;
assign COL[1106] = 1'b0;
assign COL[1107] = 1'b0;
assign COL[1108] = 1'b0;
assign COL[1109] = 1'b0;
assign COL[1110] = 1'b0;
assign COL[1111] = 1'b0;
assign COL[1112] = 1'b0;
assign COL[1113] = 1'b0;
assign COL[1114] = 1'b0;
assign COL[1115] = 1'b0;
assign COL[1116] = 1'b0;
assign COL[1117] = 1'b0;
assign COL[1118] = 1'b0;
assign COL[1119] = 1'b0;
assign COL[1120] = 1'b0;
assign COL[1121] = 1'b1;
assign COL[1122] = 1'b1;
assign COL[1123] = 1'b1;
assign COL[1124] = 1'b1;
assign COL[1125] = 1'b1;
assign COL[1126] = 1'b0;
assign COL[1127] = 1'b0;
assign COL[1128] = 1'b0;
assign COL[1129] = 1'b0;
assign COL[1130] = 1'b0;
assign COL[1131] = 1'b0;
assign COL[1132] = 1'b0;
assign COL[1133] = 1'b0;
assign COL[1134] = 1'b0;
assign COL[1135] = 1'b0;
assign COL[1136] = 1'b0;
assign COL[1137] = 1'b0;
assign COL[1138] = 1'b0;
assign COL[1139] = 1'b0;
assign COL[1140] = 1'b0;
assign COL[1141] = 1'b0;
assign COL[1142] = 1'b0;
assign COL[1143] = 1'b0;
assign COL[1144] = 1'b0;
assign COL[1145] = 1'b0;
assign COL[1146] = 1'b0;
assign COL[1147] = 1'b0;
assign COL[1148] = 1'b0;
assign COL[1149] = 1'b0;
assign COL[1150] = 1'b0;
assign COL[1151] = 1'b0;
assign COL[1152] = 1'b0;
assign COL[1153] = 1'b0;
assign COL[1154] = 1'b0;
assign COL[1155] = 1'b0;
assign COL[1156] = 1'b0;
assign COL[1157] = 1'b0;
assign COL[1158] = 1'b0;
assign COL[1159] = 1'b0;
assign COL[1160] = 1'b1;
assign COL[1161] = 1'b1;
assign COL[1162] = 1'b1;
assign COL[1163] = 1'b1;
assign COL[1164] = 1'b0;
assign COL[1165] = 1'b0;
assign COL[1166] = 1'b0;
assign COL[1167] = 1'b0;
assign COL[1168] = 1'b0;
assign COL[1169] = 1'b0;
assign COL[1170] = 1'b0;
assign COL[1171] = 1'b0;
assign COL[1172] = 1'b0;
assign COL[1173] = 1'b0;
assign COL[1174] = 1'b0;
assign COL[1175] = 1'b0;
assign COL[1176] = 1'b0;
assign COL[1177] = 1'b0;
assign COL[1178] = 1'b0;
assign COL[1179] = 1'b0;
assign COL[1180] = 1'b0;
assign COL[1181] = 1'b0;
assign COL[1182] = 1'b0;
assign COL[1183] = 1'b0;
assign COL[1184] = 1'b0;
assign COL[1185] = 1'b0;
assign COL[1186] = 1'b0;
assign COL[1187] = 1'b0;
assign COL[1188] = 1'b0;
assign COL[1189] = 1'b0;
assign COL[1190] = 1'b0;
assign COL[1191] = 1'b0;
assign COL[1192] = 1'b1;
assign COL[1193] = 1'b1;
assign COL[1194] = 1'b1;
assign COL[1195] = 1'b1;
assign COL[1196] = 1'b0;
assign COL[1197] = 1'b0;
assign COL[1198] = 1'b0;
assign COL[1199] = 1'b0;
assign COL[1200] = 1'b0;
assign COL[1201] = 1'b0;
assign COL[1202] = 1'b0;
assign COL[1203] = 1'b0;
assign COL[1204] = 1'b0;
assign COL[1205] = 1'b0;
assign COL[1206] = 1'b0;
assign COL[1207] = 1'b0;
assign COL[1208] = 1'b0;
assign COL[1209] = 1'b0;
assign COL[1210] = 1'b1;
assign COL[1211] = 1'b1;
assign COL[1212] = 1'b1;
assign COL[1213] = 1'b1;
assign COL[1214] = 1'b1;
assign COL[1215] = 1'b0;
assign COL[1216] = 1'b0;
assign COL[1217] = 1'b0;
assign COL[1218] = 1'b0;
assign COL[1219] = 1'b0;
assign COL[1220] = 1'b0;
assign COL[1221] = 1'b0;
assign COL[1222] = 1'b0;
assign COL[1223] = 1'b0;
assign COL[1224] = 1'b0;
assign COL[1225] = 1'b0;
assign COL[1226] = 1'b0;
assign COL[1227] = 1'b0;
assign COL[1228] = 1'b0;
assign COL[1229] = 1'b0;
assign COL[1230] = 1'b0;
assign COL[1231] = 1'b0;
assign COL[1232] = 1'b0;
assign COL[1233] = 1'b0;
assign COL[1234] = 1'b0;
assign COL[1235] = 1'b0;
assign COL[1236] = 1'b0;
assign COL[1237] = 1'b0;
assign COL[1238] = 1'b0;
assign COL[1239] = 1'b0;
assign COL[1240] = 1'b0;
assign COL[1241] = 1'b0;
assign COL[1242] = 1'b0;
assign COL[1243] = 1'b0;
assign COL[1244] = 1'b0;
assign COL[1245] = 1'b0;
assign COL[1246] = 1'b0;
assign COL[1247] = 1'b0;
assign COL[1248] = 1'b0;
assign COL[1249] = 1'b0;
assign COL[1250] = 1'b0;
assign COL[1251] = 1'b0;
assign COL[1252] = 1'b0;
assign COL[1253] = 1'b0;
assign COL[1254] = 1'b0;
assign COL[1255] = 1'b0;
assign COL[1256] = 1'b0;
assign COL[1257] = 1'b0;
assign COL[1258] = 1'b0;
assign COL[1259] = 1'b0;
assign COL[1260] = 1'b0;
assign COL[1261] = 1'b0;
assign COL[1262] = 1'b0;
assign COL[1263] = 1'b0;
assign COL[1264] = 1'b0;
assign COL[1265] = 1'b0;
assign COL[1266] = 1'b0;
assign COL[1267] = 1'b0;
assign COL[1268] = 1'b0;
assign COL[1269] = 1'b0;
assign COL[1270] = 1'b0;
assign COL[1271] = 1'b0;
assign COL[1272] = 1'b0;
assign COL[1273] = 1'b0;
assign COL[1274] = 1'b0;
assign COL[1275] = 1'b0;
assign COL[1276] = 1'b0;
assign COL[1277] = 1'b0;
assign COL[1278] = 1'b0;
assign COL[1279] = 1'b0;
assign COL[1280] = 1'b0;
assign COL[1281] = 1'b1;
assign COL[1282] = 1'b1;
assign COL[1283] = 1'b1;
assign COL[1284] = 1'b1;
assign COL[1285] = 1'b1;
assign COL[1286] = 1'b0;
assign COL[1287] = 1'b0;
assign COL[1288] = 1'b0;
assign COL[1289] = 1'b0;
assign COL[1290] = 1'b0;
assign COL[1291] = 1'b0;
assign COL[1292] = 1'b0;
assign COL[1293] = 1'b0;
assign COL[1294] = 1'b0;
assign COL[1295] = 1'b0;
assign COL[1296] = 1'b0;
assign COL[1297] = 1'b0;
assign COL[1298] = 1'b0;
assign COL[1299] = 1'b0;
assign COL[1300] = 1'b0;
assign COL[1301] = 1'b0;
assign COL[1302] = 1'b0;
assign COL[1303] = 1'b0;
assign COL[1304] = 1'b0;
assign COL[1305] = 1'b0;
assign COL[1306] = 1'b0;
assign COL[1307] = 1'b0;
assign COL[1308] = 1'b0;
assign COL[1309] = 1'b0;
assign COL[1310] = 1'b0;
assign COL[1311] = 1'b0;
assign COL[1312] = 1'b0;
assign COL[1313] = 1'b0;
assign COL[1314] = 1'b0;
assign COL[1315] = 1'b0;
assign COL[1316] = 1'b0;
assign COL[1317] = 1'b0;
assign COL[1318] = 1'b0;
assign COL[1319] = 1'b0;
assign COL[1320] = 1'b1;
assign COL[1321] = 1'b1;
assign COL[1322] = 1'b1;
assign COL[1323] = 1'b1;
assign COL[1324] = 1'b0;
assign COL[1325] = 1'b0;
assign COL[1326] = 1'b0;
assign COL[1327] = 1'b0;
assign COL[1328] = 1'b0;
assign COL[1329] = 1'b0;
assign COL[1330] = 1'b0;
assign COL[1331] = 1'b0;
assign COL[1332] = 1'b0;
assign COL[1333] = 1'b0;
assign COL[1334] = 1'b0;
assign COL[1335] = 1'b0;
assign COL[1336] = 1'b0;
assign COL[1337] = 1'b0;
assign COL[1338] = 1'b0;
assign COL[1339] = 1'b0;
assign COL[1340] = 1'b0;
assign COL[1341] = 1'b0;
assign COL[1342] = 1'b0;
assign COL[1343] = 1'b0;
assign COL[1344] = 1'b0;
assign COL[1345] = 1'b0;
assign COL[1346] = 1'b0;
assign COL[1347] = 1'b0;
assign COL[1348] = 1'b0;
assign COL[1349] = 1'b0;
assign COL[1350] = 1'b0;
assign COL[1351] = 1'b0;
assign COL[1352] = 1'b1;
assign COL[1353] = 1'b1;
assign COL[1354] = 1'b1;
assign COL[1355] = 1'b1;
assign COL[1356] = 1'b0;
assign COL[1357] = 1'b0;
assign COL[1358] = 1'b0;
assign COL[1359] = 1'b0;
assign COL[1360] = 1'b0;
assign COL[1361] = 1'b0;
assign COL[1362] = 1'b0;
assign COL[1363] = 1'b0;
assign COL[1364] = 1'b0;
assign COL[1365] = 1'b0;
assign COL[1366] = 1'b0;
assign COL[1367] = 1'b0;
assign COL[1368] = 1'b0;
assign COL[1369] = 1'b0;
assign COL[1370] = 1'b1;
assign COL[1371] = 1'b1;
assign COL[1372] = 1'b1;
assign COL[1373] = 1'b1;
assign COL[1374] = 1'b1;
assign COL[1375] = 1'b0;
assign COL[1376] = 1'b0;
assign COL[1377] = 1'b0;
assign COL[1378] = 1'b0;
assign COL[1379] = 1'b0;
assign COL[1380] = 1'b0;
assign COL[1381] = 1'b0;
assign COL[1382] = 1'b0;
assign COL[1383] = 1'b0;
assign COL[1384] = 1'b0;
assign COL[1385] = 1'b0;
assign COL[1386] = 1'b0;
assign COL[1387] = 1'b0;
assign COL[1388] = 1'b0;
assign COL[1389] = 1'b0;
assign COL[1390] = 1'b0;
assign COL[1391] = 1'b0;
assign COL[1392] = 1'b0;
assign COL[1393] = 1'b0;
assign COL[1394] = 1'b0;
assign COL[1395] = 1'b0;
assign COL[1396] = 1'b0;
assign COL[1397] = 1'b0;
assign COL[1398] = 1'b0;
assign COL[1399] = 1'b0;
assign COL[1400] = 1'b0;
assign COL[1401] = 1'b0;
assign COL[1402] = 1'b0;
assign COL[1403] = 1'b0;
assign COL[1404] = 1'b0;
assign COL[1405] = 1'b0;
assign COL[1406] = 1'b0;
assign COL[1407] = 1'b0;
assign COL[1408] = 1'b0;
assign COL[1409] = 1'b0;
assign COL[1410] = 1'b0;
assign COL[1411] = 1'b0;
assign COL[1412] = 1'b0;
assign COL[1413] = 1'b0;
assign COL[1414] = 1'b0;
assign COL[1415] = 1'b0;
assign COL[1416] = 1'b0;
assign COL[1417] = 1'b0;
assign COL[1418] = 1'b0;
assign COL[1419] = 1'b0;
assign COL[1420] = 1'b0;
assign COL[1421] = 1'b0;
assign COL[1422] = 1'b0;
assign COL[1423] = 1'b0;
assign COL[1424] = 1'b0;
assign COL[1425] = 1'b0;
assign COL[1426] = 1'b0;
assign COL[1427] = 1'b0;
assign COL[1428] = 1'b0;
assign COL[1429] = 1'b0;
assign COL[1430] = 1'b0;
assign COL[1431] = 1'b0;
assign COL[1432] = 1'b0;
assign COL[1433] = 1'b0;
assign COL[1434] = 1'b0;
assign COL[1435] = 1'b0;
assign COL[1436] = 1'b0;
assign COL[1437] = 1'b0;
assign COL[1438] = 1'b0;
assign COL[1439] = 1'b0;
assign COL[1440] = 1'b0;
assign COL[1441] = 1'b1;
assign COL[1442] = 1'b1;
assign COL[1443] = 1'b1;
assign COL[1444] = 1'b1;
assign COL[1445] = 1'b1;
assign COL[1446] = 1'b0;
assign COL[1447] = 1'b0;
assign COL[1448] = 1'b0;
assign COL[1449] = 1'b0;
assign COL[1450] = 1'b0;
assign COL[1451] = 1'b0;
assign COL[1452] = 1'b0;
assign COL[1453] = 1'b0;
assign COL[1454] = 1'b0;
assign COL[1455] = 1'b0;
assign COL[1456] = 1'b0;
assign COL[1457] = 1'b0;
assign COL[1458] = 1'b0;
assign COL[1459] = 1'b0;
assign COL[1460] = 1'b0;
assign COL[1461] = 1'b0;
assign COL[1462] = 1'b0;
assign COL[1463] = 1'b0;
assign COL[1464] = 1'b0;
assign COL[1465] = 1'b0;
assign COL[1466] = 1'b0;
assign COL[1467] = 1'b0;
assign COL[1468] = 1'b0;
assign COL[1469] = 1'b0;
assign COL[1470] = 1'b0;
assign COL[1471] = 1'b0;
assign COL[1472] = 1'b0;
assign COL[1473] = 1'b0;
assign COL[1474] = 1'b0;
assign COL[1475] = 1'b0;
assign COL[1476] = 1'b0;
assign COL[1477] = 1'b0;
assign COL[1478] = 1'b0;
assign COL[1479] = 1'b0;
assign COL[1480] = 1'b1;
assign COL[1481] = 1'b1;
assign COL[1482] = 1'b1;
assign COL[1483] = 1'b1;
assign COL[1484] = 1'b0;
assign COL[1485] = 1'b0;
assign COL[1486] = 1'b0;
assign COL[1487] = 1'b0;
assign COL[1488] = 1'b0;
assign COL[1489] = 1'b0;
assign COL[1490] = 1'b0;
assign COL[1491] = 1'b0;
assign COL[1492] = 1'b0;
assign COL[1493] = 1'b0;
assign COL[1494] = 1'b0;
assign COL[1495] = 1'b0;
assign COL[1496] = 1'b0;
assign COL[1497] = 1'b0;
assign COL[1498] = 1'b0;
assign COL[1499] = 1'b0;
assign COL[1500] = 1'b0;
assign COL[1501] = 1'b0;
assign COL[1502] = 1'b0;
assign COL[1503] = 1'b0;
assign COL[1504] = 1'b0;
assign COL[1505] = 1'b0;
assign COL[1506] = 1'b0;
assign COL[1507] = 1'b0;
assign COL[1508] = 1'b0;
assign COL[1509] = 1'b0;
assign COL[1510] = 1'b0;
assign COL[1511] = 1'b0;
assign COL[1512] = 1'b1;
assign COL[1513] = 1'b1;
assign COL[1514] = 1'b1;
assign COL[1515] = 1'b1;
assign COL[1516] = 1'b0;
assign COL[1517] = 1'b0;
assign COL[1518] = 1'b0;
assign COL[1519] = 1'b0;
assign COL[1520] = 1'b0;
assign COL[1521] = 1'b0;
assign COL[1522] = 1'b0;
assign COL[1523] = 1'b0;
assign COL[1524] = 1'b0;
assign COL[1525] = 1'b0;
assign COL[1526] = 1'b0;
assign COL[1527] = 1'b0;
assign COL[1528] = 1'b0;
assign COL[1529] = 1'b0;
assign COL[1530] = 1'b1;
assign COL[1531] = 1'b1;
assign COL[1532] = 1'b1;
assign COL[1533] = 1'b1;
assign COL[1534] = 1'b1;
assign COL[1535] = 1'b0;
assign COL[1536] = 1'b0;
assign COL[1537] = 1'b0;
assign COL[1538] = 1'b0;
assign COL[1539] = 1'b0;
assign COL[1540] = 1'b0;
assign COL[1541] = 1'b0;
assign COL[1542] = 1'b0;
assign COL[1543] = 1'b0;
assign COL[1544] = 1'b0;
assign COL[1545] = 1'b0;
assign COL[1546] = 1'b0;
assign COL[1547] = 1'b0;
assign COL[1548] = 1'b0;
assign COL[1549] = 1'b0;
assign COL[1550] = 1'b0;
assign COL[1551] = 1'b0;
assign COL[1552] = 1'b0;
assign COL[1553] = 1'b0;
assign COL[1554] = 1'b0;
assign COL[1555] = 1'b0;
assign COL[1556] = 1'b0;
assign COL[1557] = 1'b0;
assign COL[1558] = 1'b0;
assign COL[1559] = 1'b0;
assign COL[1560] = 1'b0;
assign COL[1561] = 1'b0;
assign COL[1562] = 1'b0;
assign COL[1563] = 1'b0;
assign COL[1564] = 1'b0;
assign COL[1565] = 1'b0;
assign COL[1566] = 1'b0;
assign COL[1567] = 1'b0;
assign COL[1568] = 1'b0;
assign COL[1569] = 1'b0;
assign COL[1570] = 1'b0;
assign COL[1571] = 1'b0;
assign COL[1572] = 1'b0;
assign COL[1573] = 1'b0;
assign COL[1574] = 1'b0;
assign COL[1575] = 1'b0;
assign COL[1576] = 1'b0;
assign COL[1577] = 1'b0;
assign COL[1578] = 1'b0;
assign COL[1579] = 1'b0;
assign COL[1580] = 1'b0;
assign COL[1581] = 1'b0;
assign COL[1582] = 1'b0;
assign COL[1583] = 1'b0;
assign COL[1584] = 1'b0;
assign COL[1585] = 1'b0;
assign COL[1586] = 1'b0;
assign COL[1587] = 1'b0;
assign COL[1588] = 1'b0;
assign COL[1589] = 1'b0;
assign COL[1590] = 1'b0;
assign COL[1591] = 1'b0;
assign COL[1592] = 1'b0;
assign COL[1593] = 1'b0;
assign COL[1594] = 1'b0;
assign COL[1595] = 1'b0;
assign COL[1596] = 1'b0;
assign COL[1597] = 1'b0;
assign COL[1598] = 1'b0;
assign COL[1599] = 1'b0;
assign COL[1600] = 1'b0;
assign COL[1601] = 1'b1;
assign COL[1602] = 1'b1;
assign COL[1603] = 1'b1;
assign COL[1604] = 1'b1;
assign COL[1605] = 1'b1;
assign COL[1606] = 1'b0;
assign COL[1607] = 1'b0;
assign COL[1608] = 1'b0;
assign COL[1609] = 1'b0;
assign COL[1610] = 1'b0;
assign COL[1611] = 1'b0;
assign COL[1612] = 1'b0;
assign COL[1613] = 1'b0;
assign COL[1614] = 1'b0;
assign COL[1615] = 1'b0;
assign COL[1616] = 1'b0;
assign COL[1617] = 1'b0;
assign COL[1618] = 1'b0;
assign COL[1619] = 1'b0;
assign COL[1620] = 1'b0;
assign COL[1621] = 1'b0;
assign COL[1622] = 1'b0;
assign COL[1623] = 1'b0;
assign COL[1624] = 1'b0;
assign COL[1625] = 1'b0;
assign COL[1626] = 1'b0;
assign COL[1627] = 1'b0;
assign COL[1628] = 1'b0;
assign COL[1629] = 1'b0;
assign COL[1630] = 1'b0;
assign COL[1631] = 1'b0;
assign COL[1632] = 1'b0;
assign COL[1633] = 1'b0;
assign COL[1634] = 1'b0;
assign COL[1635] = 1'b0;
assign COL[1636] = 1'b0;
assign COL[1637] = 1'b0;
assign COL[1638] = 1'b0;
assign COL[1639] = 1'b0;
assign COL[1640] = 1'b1;
assign COL[1641] = 1'b1;
assign COL[1642] = 1'b1;
assign COL[1643] = 1'b1;
assign COL[1644] = 1'b0;
assign COL[1645] = 1'b0;
assign COL[1646] = 1'b0;
assign COL[1647] = 1'b0;
assign COL[1648] = 1'b0;
assign COL[1649] = 1'b0;
assign COL[1650] = 1'b0;
assign COL[1651] = 1'b0;
assign COL[1652] = 1'b0;
assign COL[1653] = 1'b0;
assign COL[1654] = 1'b0;
assign COL[1655] = 1'b0;
assign COL[1656] = 1'b0;
assign COL[1657] = 1'b0;
assign COL[1658] = 1'b0;
assign COL[1659] = 1'b0;
assign COL[1660] = 1'b0;
assign COL[1661] = 1'b0;
assign COL[1662] = 1'b0;
assign COL[1663] = 1'b0;
assign COL[1664] = 1'b0;
assign COL[1665] = 1'b0;
assign COL[1666] = 1'b0;
assign COL[1667] = 1'b0;
assign COL[1668] = 1'b0;
assign COL[1669] = 1'b0;
assign COL[1670] = 1'b0;
assign COL[1671] = 1'b0;
assign COL[1672] = 1'b1;
assign COL[1673] = 1'b1;
assign COL[1674] = 1'b1;
assign COL[1675] = 1'b1;
assign COL[1676] = 1'b0;
assign COL[1677] = 1'b0;
assign COL[1678] = 1'b0;
assign COL[1679] = 1'b0;
assign COL[1680] = 1'b0;
assign COL[1681] = 1'b0;
assign COL[1682] = 1'b0;
assign COL[1683] = 1'b0;
assign COL[1684] = 1'b0;
assign COL[1685] = 1'b0;
assign COL[1686] = 1'b0;
assign COL[1687] = 1'b0;
assign COL[1688] = 1'b0;
assign COL[1689] = 1'b0;
assign COL[1690] = 1'b1;
assign COL[1691] = 1'b1;
assign COL[1692] = 1'b1;
assign COL[1693] = 1'b1;
assign COL[1694] = 1'b1;
assign COL[1695] = 1'b0;
assign COL[1696] = 1'b0;
assign COL[1697] = 1'b0;
assign COL[1698] = 1'b0;
assign COL[1699] = 1'b0;
assign COL[1700] = 1'b0;
assign COL[1701] = 1'b0;
assign COL[1702] = 1'b0;
assign COL[1703] = 1'b0;
assign COL[1704] = 1'b0;
assign COL[1705] = 1'b0;
assign COL[1706] = 1'b0;
assign COL[1707] = 1'b0;
assign COL[1708] = 1'b0;
assign COL[1709] = 1'b0;
assign COL[1710] = 1'b0;
assign COL[1711] = 1'b0;
assign COL[1712] = 1'b0;
assign COL[1713] = 1'b0;
assign COL[1714] = 1'b0;
assign COL[1715] = 1'b0;
assign COL[1716] = 1'b0;
assign COL[1717] = 1'b0;
assign COL[1718] = 1'b0;
assign COL[1719] = 1'b0;
assign COL[1720] = 1'b0;
assign COL[1721] = 1'b0;
assign COL[1722] = 1'b0;
assign COL[1723] = 1'b0;
assign COL[1724] = 1'b0;
assign COL[1725] = 1'b0;
assign COL[1726] = 1'b0;
assign COL[1727] = 1'b0;
assign COL[1728] = 1'b0;
assign COL[1729] = 1'b0;
assign COL[1730] = 1'b0;
assign COL[1731] = 1'b0;
assign COL[1732] = 1'b0;
assign COL[1733] = 1'b0;
assign COL[1734] = 1'b0;
assign COL[1735] = 1'b0;
assign COL[1736] = 1'b0;
assign COL[1737] = 1'b0;
assign COL[1738] = 1'b0;
assign COL[1739] = 1'b0;
assign COL[1740] = 1'b0;
assign COL[1741] = 1'b0;
assign COL[1742] = 1'b0;
assign COL[1743] = 1'b0;
assign COL[1744] = 1'b0;
assign COL[1745] = 1'b0;
assign COL[1746] = 1'b0;
assign COL[1747] = 1'b0;
assign COL[1748] = 1'b0;
assign COL[1749] = 1'b0;
assign COL[1750] = 1'b0;
assign COL[1751] = 1'b0;
assign COL[1752] = 1'b0;
assign COL[1753] = 1'b0;
assign COL[1754] = 1'b0;
assign COL[1755] = 1'b0;
assign COL[1756] = 1'b0;
assign COL[1757] = 1'b0;
assign COL[1758] = 1'b0;
assign COL[1759] = 1'b0;
assign COL[1760] = 1'b0;
assign COL[1761] = 1'b1;
assign COL[1762] = 1'b1;
assign COL[1763] = 1'b1;
assign COL[1764] = 1'b1;
assign COL[1765] = 1'b1;
assign COL[1766] = 1'b0;
assign COL[1767] = 1'b0;
assign COL[1768] = 1'b0;
assign COL[1769] = 1'b0;
assign COL[1770] = 1'b0;
assign COL[1771] = 1'b0;
assign COL[1772] = 1'b0;
assign COL[1773] = 1'b0;
assign COL[1774] = 1'b0;
assign COL[1775] = 1'b0;
assign COL[1776] = 1'b0;
assign COL[1777] = 1'b0;
assign COL[1778] = 1'b0;
assign COL[1779] = 1'b0;
assign COL[1780] = 1'b0;
assign COL[1781] = 1'b0;
assign COL[1782] = 1'b0;
assign COL[1783] = 1'b0;
assign COL[1784] = 1'b0;
assign COL[1785] = 1'b0;
assign COL[1786] = 1'b0;
assign COL[1787] = 1'b0;
assign COL[1788] = 1'b0;
assign COL[1789] = 1'b0;
assign COL[1790] = 1'b0;
assign COL[1791] = 1'b0;
assign COL[1792] = 1'b0;
assign COL[1793] = 1'b0;
assign COL[1794] = 1'b0;
assign COL[1795] = 1'b0;
assign COL[1796] = 1'b0;
assign COL[1797] = 1'b0;
assign COL[1798] = 1'b0;
assign COL[1799] = 1'b0;
assign COL[1800] = 1'b1;
assign COL[1801] = 1'b1;
assign COL[1802] = 1'b1;
assign COL[1803] = 1'b1;
assign COL[1804] = 1'b0;
assign COL[1805] = 1'b0;
assign COL[1806] = 1'b0;
assign COL[1807] = 1'b0;
assign COL[1808] = 1'b0;
assign COL[1809] = 1'b0;
assign COL[1810] = 1'b0;
assign COL[1811] = 1'b0;
assign COL[1812] = 1'b0;
assign COL[1813] = 1'b0;
assign COL[1814] = 1'b0;
assign COL[1815] = 1'b0;
assign COL[1816] = 1'b0;
assign COL[1817] = 1'b0;
assign COL[1818] = 1'b0;
assign COL[1819] = 1'b0;
assign COL[1820] = 1'b0;
assign COL[1821] = 1'b0;
assign COL[1822] = 1'b0;
assign COL[1823] = 1'b0;
assign COL[1824] = 1'b0;
assign COL[1825] = 1'b0;
assign COL[1826] = 1'b0;
assign COL[1827] = 1'b0;
assign COL[1828] = 1'b0;
assign COL[1829] = 1'b0;
assign COL[1830] = 1'b0;
assign COL[1831] = 1'b0;
assign COL[1832] = 1'b1;
assign COL[1833] = 1'b1;
assign COL[1834] = 1'b1;
assign COL[1835] = 1'b1;
assign COL[1836] = 1'b0;
assign COL[1837] = 1'b0;
assign COL[1838] = 1'b0;
assign COL[1839] = 1'b0;
assign COL[1840] = 1'b0;
assign COL[1841] = 1'b0;
assign COL[1842] = 1'b0;
assign COL[1843] = 1'b0;
assign COL[1844] = 1'b0;
assign COL[1845] = 1'b0;
assign COL[1846] = 1'b0;
assign COL[1847] = 1'b0;
assign COL[1848] = 1'b0;
assign COL[1849] = 1'b0;
assign COL[1850] = 1'b1;
assign COL[1851] = 1'b1;
assign COL[1852] = 1'b1;
assign COL[1853] = 1'b1;
assign COL[1854] = 1'b1;
assign COL[1855] = 1'b0;
assign COL[1856] = 1'b0;
assign COL[1857] = 1'b0;
assign COL[1858] = 1'b0;
assign COL[1859] = 1'b0;
assign COL[1860] = 1'b0;
assign COL[1861] = 1'b0;
assign COL[1862] = 1'b0;
assign COL[1863] = 1'b0;
assign COL[1864] = 1'b0;
assign COL[1865] = 1'b0;
assign COL[1866] = 1'b0;
assign COL[1867] = 1'b0;
assign COL[1868] = 1'b0;
assign COL[1869] = 1'b0;
assign COL[1870] = 1'b0;
assign COL[1871] = 1'b0;
assign COL[1872] = 1'b0;
assign COL[1873] = 1'b0;
assign COL[1874] = 1'b0;
assign COL[1875] = 1'b0;
assign COL[1876] = 1'b0;
assign COL[1877] = 1'b0;
assign COL[1878] = 1'b0;
assign COL[1879] = 1'b0;
assign COL[1880] = 1'b0;
assign COL[1881] = 1'b0;
assign COL[1882] = 1'b0;
assign COL[1883] = 1'b0;
assign COL[1884] = 1'b0;
assign COL[1885] = 1'b0;
assign COL[1886] = 1'b0;
assign COL[1887] = 1'b0;
assign COL[1888] = 1'b0;
assign COL[1889] = 1'b0;
assign COL[1890] = 1'b0;
assign COL[1891] = 1'b0;
assign COL[1892] = 1'b0;
assign COL[1893] = 1'b0;
assign COL[1894] = 1'b0;
assign COL[1895] = 1'b0;
assign COL[1896] = 1'b0;
assign COL[1897] = 1'b0;
assign COL[1898] = 1'b0;
assign COL[1899] = 1'b0;
assign COL[1900] = 1'b0;
assign COL[1901] = 1'b0;
assign COL[1902] = 1'b0;
assign COL[1903] = 1'b0;
assign COL[1904] = 1'b0;
assign COL[1905] = 1'b0;
assign COL[1906] = 1'b0;
assign COL[1907] = 1'b0;
assign COL[1908] = 1'b0;
assign COL[1909] = 1'b0;
assign COL[1910] = 1'b0;
assign COL[1911] = 1'b0;
assign COL[1912] = 1'b0;
assign COL[1913] = 1'b0;
assign COL[1914] = 1'b0;
assign COL[1915] = 1'b0;
assign COL[1916] = 1'b0;
assign COL[1917] = 1'b0;
assign COL[1918] = 1'b0;
assign COL[1919] = 1'b0;
assign COL[1920] = 1'b0;
assign COL[1921] = 1'b1;
assign COL[1922] = 1'b1;
assign COL[1923] = 1'b1;
assign COL[1924] = 1'b1;
assign COL[1925] = 1'b1;
assign COL[1926] = 1'b0;
assign COL[1927] = 1'b0;
assign COL[1928] = 1'b0;
assign COL[1929] = 1'b0;
assign COL[1930] = 1'b0;
assign COL[1931] = 1'b0;
assign COL[1932] = 1'b0;
assign COL[1933] = 1'b0;
assign COL[1934] = 1'b0;
assign COL[1935] = 1'b0;
assign COL[1936] = 1'b0;
assign COL[1937] = 1'b0;
assign COL[1938] = 1'b0;
assign COL[1939] = 1'b0;
assign COL[1940] = 1'b0;
assign COL[1941] = 1'b0;
assign COL[1942] = 1'b0;
assign COL[1943] = 1'b0;
assign COL[1944] = 1'b0;
assign COL[1945] = 1'b0;
assign COL[1946] = 1'b0;
assign COL[1947] = 1'b0;
assign COL[1948] = 1'b0;
assign COL[1949] = 1'b0;
assign COL[1950] = 1'b0;
assign COL[1951] = 1'b0;
assign COL[1952] = 1'b0;
assign COL[1953] = 1'b0;
assign COL[1954] = 1'b0;
assign COL[1955] = 1'b0;
assign COL[1956] = 1'b0;
assign COL[1957] = 1'b0;
assign COL[1958] = 1'b0;
assign COL[1959] = 1'b0;
assign COL[1960] = 1'b1;
assign COL[1961] = 1'b1;
assign COL[1962] = 1'b1;
assign COL[1963] = 1'b1;
assign COL[1964] = 1'b0;
assign COL[1965] = 1'b0;
assign COL[1966] = 1'b0;
assign COL[1967] = 1'b0;
assign COL[1968] = 1'b0;
assign COL[1969] = 1'b0;
assign COL[1970] = 1'b0;
assign COL[1971] = 1'b0;
assign COL[1972] = 1'b0;
assign COL[1973] = 1'b0;
assign COL[1974] = 1'b0;
assign COL[1975] = 1'b0;
assign COL[1976] = 1'b0;
assign COL[1977] = 1'b0;
assign COL[1978] = 1'b0;
assign COL[1979] = 1'b0;
assign COL[1980] = 1'b0;
assign COL[1981] = 1'b0;
assign COL[1982] = 1'b0;
assign COL[1983] = 1'b0;
assign COL[1984] = 1'b0;
assign COL[1985] = 1'b0;
assign COL[1986] = 1'b0;
assign COL[1987] = 1'b0;
assign COL[1988] = 1'b0;
assign COL[1989] = 1'b0;
assign COL[1990] = 1'b0;
assign COL[1991] = 1'b0;
assign COL[1992] = 1'b1;
assign COL[1993] = 1'b1;
assign COL[1994] = 1'b1;
assign COL[1995] = 1'b1;
assign COL[1996] = 1'b0;
assign COL[1997] = 1'b0;
assign COL[1998] = 1'b0;
assign COL[1999] = 1'b0;
assign COL[2000] = 1'b0;
assign COL[2001] = 1'b0;
assign COL[2002] = 1'b0;
assign COL[2003] = 1'b0;
assign COL[2004] = 1'b0;
assign COL[2005] = 1'b0;
assign COL[2006] = 1'b0;
assign COL[2007] = 1'b0;
assign COL[2008] = 1'b0;
assign COL[2009] = 1'b0;
assign COL[2010] = 1'b1;
assign COL[2011] = 1'b1;
assign COL[2012] = 1'b1;
assign COL[2013] = 1'b1;
assign COL[2014] = 1'b1;
assign COL[2015] = 1'b0;
assign COL[2016] = 1'b0;
assign COL[2017] = 1'b0;
assign COL[2018] = 1'b0;
assign COL[2019] = 1'b0;
assign COL[2020] = 1'b0;
assign COL[2021] = 1'b0;
assign COL[2022] = 1'b0;
assign COL[2023] = 1'b0;
assign COL[2024] = 1'b0;
assign COL[2025] = 1'b0;
assign COL[2026] = 1'b0;
assign COL[2027] = 1'b0;
assign COL[2028] = 1'b0;
assign COL[2029] = 1'b0;
assign COL[2030] = 1'b0;
assign COL[2031] = 1'b0;
assign COL[2032] = 1'b0;
assign COL[2033] = 1'b0;
assign COL[2034] = 1'b0;
assign COL[2035] = 1'b0;
assign COL[2036] = 1'b0;
assign COL[2037] = 1'b0;
assign COL[2038] = 1'b0;
assign COL[2039] = 1'b0;
assign COL[2040] = 1'b0;
assign COL[2041] = 1'b0;
assign COL[2042] = 1'b0;
assign COL[2043] = 1'b0;
assign COL[2044] = 1'b0;
assign COL[2045] = 1'b0;
assign COL[2046] = 1'b0;
assign COL[2047] = 1'b0;
assign COL[2048] = 1'b0;
assign COL[2049] = 1'b0;
assign COL[2050] = 1'b0;
assign COL[2051] = 1'b0;
assign COL[2052] = 1'b0;
assign COL[2053] = 1'b0;
assign COL[2054] = 1'b0;
assign COL[2055] = 1'b0;
assign COL[2056] = 1'b0;
assign COL[2057] = 1'b0;
assign COL[2058] = 1'b0;
assign COL[2059] = 1'b0;
assign COL[2060] = 1'b0;
assign COL[2061] = 1'b0;
assign COL[2062] = 1'b0;
assign COL[2063] = 1'b0;
assign COL[2064] = 1'b0;
assign COL[2065] = 1'b0;
assign COL[2066] = 1'b0;
assign COL[2067] = 1'b0;
assign COL[2068] = 1'b0;
assign COL[2069] = 1'b0;
assign COL[2070] = 1'b0;
assign COL[2071] = 1'b0;
assign COL[2072] = 1'b0;
assign COL[2073] = 1'b0;
assign COL[2074] = 1'b0;
assign COL[2075] = 1'b0;
assign COL[2076] = 1'b0;
assign COL[2077] = 1'b0;
assign COL[2078] = 1'b0;
assign COL[2079] = 1'b0;
assign COL[2080] = 1'b0;
assign COL[2081] = 1'b1;
assign COL[2082] = 1'b1;
assign COL[2083] = 1'b1;
assign COL[2084] = 1'b1;
assign COL[2085] = 1'b1;
assign COL[2086] = 1'b0;
assign COL[2087] = 1'b0;
assign COL[2088] = 1'b0;
assign COL[2089] = 1'b0;
assign COL[2090] = 1'b0;
assign COL[2091] = 1'b0;
assign COL[2092] = 1'b0;
assign COL[2093] = 1'b0;
assign COL[2094] = 1'b0;
assign COL[2095] = 1'b0;
assign COL[2096] = 1'b0;
assign COL[2097] = 1'b0;
assign COL[2098] = 1'b0;
assign COL[2099] = 1'b0;
assign COL[2100] = 1'b0;
assign COL[2101] = 1'b0;
assign COL[2102] = 1'b0;
assign COL[2103] = 1'b0;
assign COL[2104] = 1'b0;
assign COL[2105] = 1'b0;
assign COL[2106] = 1'b0;
assign COL[2107] = 1'b0;
assign COL[2108] = 1'b0;
assign COL[2109] = 1'b0;
assign COL[2110] = 1'b0;
assign COL[2111] = 1'b0;
assign COL[2112] = 1'b0;
assign COL[2113] = 1'b0;
assign COL[2114] = 1'b0;
assign COL[2115] = 1'b0;
assign COL[2116] = 1'b0;
assign COL[2117] = 1'b0;
assign COL[2118] = 1'b0;
assign COL[2119] = 1'b0;
assign COL[2120] = 1'b1;
assign COL[2121] = 1'b1;
assign COL[2122] = 1'b1;
assign COL[2123] = 1'b1;
assign COL[2124] = 1'b0;
assign COL[2125] = 1'b0;
assign COL[2126] = 1'b0;
assign COL[2127] = 1'b0;
assign COL[2128] = 1'b0;
assign COL[2129] = 1'b0;
assign COL[2130] = 1'b0;
assign COL[2131] = 1'b0;
assign COL[2132] = 1'b0;
assign COL[2133] = 1'b0;
assign COL[2134] = 1'b0;
assign COL[2135] = 1'b0;
assign COL[2136] = 1'b0;
assign COL[2137] = 1'b0;
assign COL[2138] = 1'b0;
assign COL[2139] = 1'b0;
assign COL[2140] = 1'b0;
assign COL[2141] = 1'b0;
assign COL[2142] = 1'b0;
assign COL[2143] = 1'b0;
assign COL[2144] = 1'b0;
assign COL[2145] = 1'b0;
assign COL[2146] = 1'b0;
assign COL[2147] = 1'b0;
assign COL[2148] = 1'b0;
assign COL[2149] = 1'b0;
assign COL[2150] = 1'b0;
assign COL[2151] = 1'b0;
assign COL[2152] = 1'b1;
assign COL[2153] = 1'b1;
assign COL[2154] = 1'b1;
assign COL[2155] = 1'b1;
assign COL[2156] = 1'b0;
assign COL[2157] = 1'b0;
assign COL[2158] = 1'b0;
assign COL[2159] = 1'b0;
assign COL[2160] = 1'b0;
assign COL[2161] = 1'b0;
assign COL[2162] = 1'b0;
assign COL[2163] = 1'b0;
assign COL[2164] = 1'b0;
assign COL[2165] = 1'b0;
assign COL[2166] = 1'b0;
assign COL[2167] = 1'b0;
assign COL[2168] = 1'b0;
assign COL[2169] = 1'b0;
assign COL[2170] = 1'b1;
assign COL[2171] = 1'b1;
assign COL[2172] = 1'b1;
assign COL[2173] = 1'b1;
assign COL[2174] = 1'b1;
assign COL[2175] = 1'b0;
assign COL[2176] = 1'b0;
assign COL[2177] = 1'b0;
assign COL[2178] = 1'b0;
assign COL[2179] = 1'b0;
assign COL[2180] = 1'b0;
assign COL[2181] = 1'b0;
assign COL[2182] = 1'b0;
assign COL[2183] = 1'b0;
assign COL[2184] = 1'b0;
assign COL[2185] = 1'b0;
assign COL[2186] = 1'b0;
assign COL[2187] = 1'b0;
assign COL[2188] = 1'b0;
assign COL[2189] = 1'b0;
assign COL[2190] = 1'b0;
assign COL[2191] = 1'b0;
assign COL[2192] = 1'b0;
assign COL[2193] = 1'b0;
assign COL[2194] = 1'b0;
assign COL[2195] = 1'b0;
assign COL[2196] = 1'b0;
assign COL[2197] = 1'b0;
assign COL[2198] = 1'b0;
assign COL[2199] = 1'b0;
assign COL[2200] = 1'b0;
assign COL[2201] = 1'b0;
assign COL[2202] = 1'b0;
assign COL[2203] = 1'b0;
assign COL[2204] = 1'b0;
assign COL[2205] = 1'b0;
assign COL[2206] = 1'b0;
assign COL[2207] = 1'b0;
assign COL[2208] = 1'b0;
assign COL[2209] = 1'b0;
assign COL[2210] = 1'b0;
assign COL[2211] = 1'b0;
assign COL[2212] = 1'b0;
assign COL[2213] = 1'b0;
assign COL[2214] = 1'b0;
assign COL[2215] = 1'b0;
assign COL[2216] = 1'b0;
assign COL[2217] = 1'b0;
assign COL[2218] = 1'b0;
assign COL[2219] = 1'b0;
assign COL[2220] = 1'b0;
assign COL[2221] = 1'b0;
assign COL[2222] = 1'b0;
assign COL[2223] = 1'b0;
assign COL[2224] = 1'b0;
assign COL[2225] = 1'b0;
assign COL[2226] = 1'b0;
assign COL[2227] = 1'b0;
assign COL[2228] = 1'b0;
assign COL[2229] = 1'b0;
assign COL[2230] = 1'b0;
assign COL[2231] = 1'b0;
assign COL[2232] = 1'b0;
assign COL[2233] = 1'b0;
assign COL[2234] = 1'b0;
assign COL[2235] = 1'b0;
assign COL[2236] = 1'b0;
assign COL[2237] = 1'b0;
assign COL[2238] = 1'b0;
assign COL[2239] = 1'b0;
assign COL[2240] = 1'b0;
assign COL[2241] = 1'b1;
assign COL[2242] = 1'b1;
assign COL[2243] = 1'b1;
assign COL[2244] = 1'b1;
assign COL[2245] = 1'b1;
assign COL[2246] = 1'b0;
assign COL[2247] = 1'b0;
assign COL[2248] = 1'b0;
assign COL[2249] = 1'b0;
assign COL[2250] = 1'b0;
assign COL[2251] = 1'b0;
assign COL[2252] = 1'b0;
assign COL[2253] = 1'b0;
assign COL[2254] = 1'b0;
assign COL[2255] = 1'b0;
assign COL[2256] = 1'b0;
assign COL[2257] = 1'b0;
assign COL[2258] = 1'b0;
assign COL[2259] = 1'b0;
assign COL[2260] = 1'b0;
assign COL[2261] = 1'b0;
assign COL[2262] = 1'b0;
assign COL[2263] = 1'b0;
assign COL[2264] = 1'b0;
assign COL[2265] = 1'b0;
assign COL[2266] = 1'b0;
assign COL[2267] = 1'b0;
assign COL[2268] = 1'b0;
assign COL[2269] = 1'b0;
assign COL[2270] = 1'b0;
assign COL[2271] = 1'b0;
assign COL[2272] = 1'b0;
assign COL[2273] = 1'b0;
assign COL[2274] = 1'b0;
assign COL[2275] = 1'b0;
assign COL[2276] = 1'b0;
assign COL[2277] = 1'b0;
assign COL[2278] = 1'b0;
assign COL[2279] = 1'b0;
assign COL[2280] = 1'b1;
assign COL[2281] = 1'b1;
assign COL[2282] = 1'b1;
assign COL[2283] = 1'b1;
assign COL[2284] = 1'b0;
assign COL[2285] = 1'b0;
assign COL[2286] = 1'b0;
assign COL[2287] = 1'b0;
assign COL[2288] = 1'b0;
assign COL[2289] = 1'b0;
assign COL[2290] = 1'b0;
assign COL[2291] = 1'b0;
assign COL[2292] = 1'b0;
assign COL[2293] = 1'b0;
assign COL[2294] = 1'b0;
assign COL[2295] = 1'b0;
assign COL[2296] = 1'b0;
assign COL[2297] = 1'b0;
assign COL[2298] = 1'b0;
assign COL[2299] = 1'b0;
assign COL[2300] = 1'b0;
assign COL[2301] = 1'b0;
assign COL[2302] = 1'b0;
assign COL[2303] = 1'b0;
assign COL[2304] = 1'b0;
assign COL[2305] = 1'b0;
assign COL[2306] = 1'b0;
assign COL[2307] = 1'b0;
assign COL[2308] = 1'b0;
assign COL[2309] = 1'b0;
assign COL[2310] = 1'b0;
assign COL[2311] = 1'b0;
assign COL[2312] = 1'b1;
assign COL[2313] = 1'b1;
assign COL[2314] = 1'b1;
assign COL[2315] = 1'b1;
assign COL[2316] = 1'b0;
assign COL[2317] = 1'b0;
assign COL[2318] = 1'b0;
assign COL[2319] = 1'b0;
assign COL[2320] = 1'b0;
assign COL[2321] = 1'b0;
assign COL[2322] = 1'b0;
assign COL[2323] = 1'b0;
assign COL[2324] = 1'b0;
assign COL[2325] = 1'b0;
assign COL[2326] = 1'b0;
assign COL[2327] = 1'b0;
assign COL[2328] = 1'b0;
assign COL[2329] = 1'b0;
assign COL[2330] = 1'b1;
assign COL[2331] = 1'b1;
assign COL[2332] = 1'b1;
assign COL[2333] = 1'b1;
assign COL[2334] = 1'b1;
assign COL[2335] = 1'b0;
assign COL[2336] = 1'b0;
assign COL[2337] = 1'b0;
assign COL[2338] = 1'b0;
assign COL[2339] = 1'b0;
assign COL[2340] = 1'b0;
assign COL[2341] = 1'b0;
assign COL[2342] = 1'b0;
assign COL[2343] = 1'b0;
assign COL[2344] = 1'b0;
assign COL[2345] = 1'b0;
assign COL[2346] = 1'b0;
assign COL[2347] = 1'b0;
assign COL[2348] = 1'b0;
assign COL[2349] = 1'b0;
assign COL[2350] = 1'b0;
assign COL[2351] = 1'b0;
assign COL[2352] = 1'b0;
assign COL[2353] = 1'b0;
assign COL[2354] = 1'b0;
assign COL[2355] = 1'b0;
assign COL[2356] = 1'b0;
assign COL[2357] = 1'b0;
assign COL[2358] = 1'b0;
assign COL[2359] = 1'b0;
assign COL[2360] = 1'b0;
assign COL[2361] = 1'b0;
assign COL[2362] = 1'b0;
assign COL[2363] = 1'b0;
assign COL[2364] = 1'b0;
assign COL[2365] = 1'b0;
assign COL[2366] = 1'b0;
assign COL[2367] = 1'b0;
assign COL[2368] = 1'b0;
assign COL[2369] = 1'b0;
assign COL[2370] = 1'b0;
assign COL[2371] = 1'b0;
assign COL[2372] = 1'b0;
assign COL[2373] = 1'b0;
assign COL[2374] = 1'b0;
assign COL[2375] = 1'b0;
assign COL[2376] = 1'b0;
assign COL[2377] = 1'b0;
assign COL[2378] = 1'b0;
assign COL[2379] = 1'b0;
assign COL[2380] = 1'b0;
assign COL[2381] = 1'b0;
assign COL[2382] = 1'b0;
assign COL[2383] = 1'b0;
assign COL[2384] = 1'b0;
assign COL[2385] = 1'b0;
assign COL[2386] = 1'b0;
assign COL[2387] = 1'b0;
assign COL[2388] = 1'b0;
assign COL[2389] = 1'b0;
assign COL[2390] = 1'b0;
assign COL[2391] = 1'b0;
assign COL[2392] = 1'b0;
assign COL[2393] = 1'b0;
assign COL[2394] = 1'b0;
assign COL[2395] = 1'b0;
assign COL[2396] = 1'b0;
assign COL[2397] = 1'b0;
assign COL[2398] = 1'b0;
assign COL[2399] = 1'b0;
assign COL[2400] = 1'b0;
assign COL[2401] = 1'b1;
assign COL[2402] = 1'b1;
assign COL[2403] = 1'b1;
assign COL[2404] = 1'b1;
assign COL[2405] = 1'b1;
assign COL[2406] = 1'b0;
assign COL[2407] = 1'b0;
assign COL[2408] = 1'b0;
assign COL[2409] = 1'b0;
assign COL[2410] = 1'b0;
assign COL[2411] = 1'b0;
assign COL[2412] = 1'b0;
assign COL[2413] = 1'b0;
assign COL[2414] = 1'b0;
assign COL[2415] = 1'b0;
assign COL[2416] = 1'b0;
assign COL[2417] = 1'b0;
assign COL[2418] = 1'b0;
assign COL[2419] = 1'b0;
assign COL[2420] = 1'b0;
assign COL[2421] = 1'b0;
assign COL[2422] = 1'b0;
assign COL[2423] = 1'b0;
assign COL[2424] = 1'b0;
assign COL[2425] = 1'b0;
assign COL[2426] = 1'b0;
assign COL[2427] = 1'b0;
assign COL[2428] = 1'b0;
assign COL[2429] = 1'b0;
assign COL[2430] = 1'b0;
assign COL[2431] = 1'b0;
assign COL[2432] = 1'b0;
assign COL[2433] = 1'b0;
assign COL[2434] = 1'b0;
assign COL[2435] = 1'b0;
assign COL[2436] = 1'b0;
assign COL[2437] = 1'b0;
assign COL[2438] = 1'b0;
assign COL[2439] = 1'b0;
assign COL[2440] = 1'b1;
assign COL[2441] = 1'b1;
assign COL[2442] = 1'b1;
assign COL[2443] = 1'b1;
assign COL[2444] = 1'b0;
assign COL[2445] = 1'b0;
assign COL[2446] = 1'b0;
assign COL[2447] = 1'b0;
assign COL[2448] = 1'b0;
assign COL[2449] = 1'b0;
assign COL[2450] = 1'b0;
assign COL[2451] = 1'b0;
assign COL[2452] = 1'b0;
assign COL[2453] = 1'b0;
assign COL[2454] = 1'b0;
assign COL[2455] = 1'b0;
assign COL[2456] = 1'b0;
assign COL[2457] = 1'b0;
assign COL[2458] = 1'b0;
assign COL[2459] = 1'b0;
assign COL[2460] = 1'b0;
assign COL[2461] = 1'b0;
assign COL[2462] = 1'b0;
assign COL[2463] = 1'b0;
assign COL[2464] = 1'b0;
assign COL[2465] = 1'b0;
assign COL[2466] = 1'b0;
assign COL[2467] = 1'b0;
assign COL[2468] = 1'b0;
assign COL[2469] = 1'b0;
assign COL[2470] = 1'b0;
assign COL[2471] = 1'b0;
assign COL[2472] = 1'b1;
assign COL[2473] = 1'b1;
assign COL[2474] = 1'b1;
assign COL[2475] = 1'b1;
assign COL[2476] = 1'b0;
assign COL[2477] = 1'b0;
assign COL[2478] = 1'b0;
assign COL[2479] = 1'b0;
assign COL[2480] = 1'b0;
assign COL[2481] = 1'b0;
assign COL[2482] = 1'b0;
assign COL[2483] = 1'b0;
assign COL[2484] = 1'b0;
assign COL[2485] = 1'b0;
assign COL[2486] = 1'b0;
assign COL[2487] = 1'b0;
assign COL[2488] = 1'b0;
assign COL[2489] = 1'b0;
assign COL[2490] = 1'b1;
assign COL[2491] = 1'b1;
assign COL[2492] = 1'b1;
assign COL[2493] = 1'b1;
assign COL[2494] = 1'b1;
assign COL[2495] = 1'b0;
assign COL[2496] = 1'b0;
assign COL[2497] = 1'b0;
assign COL[2498] = 1'b0;
assign COL[2499] = 1'b0;
assign COL[2500] = 1'b0;
assign COL[2501] = 1'b0;
assign COL[2502] = 1'b0;
assign COL[2503] = 1'b0;
assign COL[2504] = 1'b0;
assign COL[2505] = 1'b0;
assign COL[2506] = 1'b0;
assign COL[2507] = 1'b0;
assign COL[2508] = 1'b0;
assign COL[2509] = 1'b0;
assign COL[2510] = 1'b0;
assign COL[2511] = 1'b0;
assign COL[2512] = 1'b0;
assign COL[2513] = 1'b0;
assign COL[2514] = 1'b0;
assign COL[2515] = 1'b0;
assign COL[2516] = 1'b0;
assign COL[2517] = 1'b0;
assign COL[2518] = 1'b0;
assign COL[2519] = 1'b0;
assign COL[2520] = 1'b0;
assign COL[2521] = 1'b0;
assign COL[2522] = 1'b0;
assign COL[2523] = 1'b0;
assign COL[2524] = 1'b0;
assign COL[2525] = 1'b0;
assign COL[2526] = 1'b0;
assign COL[2527] = 1'b0;
assign COL[2528] = 1'b0;
assign COL[2529] = 1'b0;
assign COL[2530] = 1'b0;
assign COL[2531] = 1'b0;
assign COL[2532] = 1'b0;
assign COL[2533] = 1'b0;
assign COL[2534] = 1'b0;
assign COL[2535] = 1'b0;
assign COL[2536] = 1'b0;
assign COL[2537] = 1'b0;
assign COL[2538] = 1'b0;
assign COL[2539] = 1'b0;
assign COL[2540] = 1'b0;
assign COL[2541] = 1'b0;
assign COL[2542] = 1'b0;
assign COL[2543] = 1'b0;
assign COL[2544] = 1'b0;
assign COL[2545] = 1'b0;
assign COL[2546] = 1'b0;
assign COL[2547] = 1'b0;
assign COL[2548] = 1'b0;
assign COL[2549] = 1'b0;
assign COL[2550] = 1'b0;
assign COL[2551] = 1'b0;
assign COL[2552] = 1'b0;
assign COL[2553] = 1'b0;
assign COL[2554] = 1'b0;
assign COL[2555] = 1'b0;
assign COL[2556] = 1'b0;
assign COL[2557] = 1'b0;
assign COL[2558] = 1'b0;
assign COL[2559] = 1'b0;
assign COL[2560] = 1'b0;
assign COL[2561] = 1'b1;
assign COL[2562] = 1'b1;
assign COL[2563] = 1'b1;
assign COL[2564] = 1'b1;
assign COL[2565] = 1'b1;
assign COL[2566] = 1'b0;
assign COL[2567] = 1'b0;
assign COL[2568] = 1'b0;
assign COL[2569] = 1'b0;
assign COL[2570] = 1'b0;
assign COL[2571] = 1'b0;
assign COL[2572] = 1'b0;
assign COL[2573] = 1'b0;
assign COL[2574] = 1'b0;
assign COL[2575] = 1'b0;
assign COL[2576] = 1'b0;
assign COL[2577] = 1'b0;
assign COL[2578] = 1'b0;
assign COL[2579] = 1'b0;
assign COL[2580] = 1'b0;
assign COL[2581] = 1'b0;
assign COL[2582] = 1'b0;
assign COL[2583] = 1'b0;
assign COL[2584] = 1'b0;
assign COL[2585] = 1'b0;
assign COL[2586] = 1'b0;
assign COL[2587] = 1'b0;
assign COL[2588] = 1'b0;
assign COL[2589] = 1'b0;
assign COL[2590] = 1'b0;
assign COL[2591] = 1'b0;
assign COL[2592] = 1'b0;
assign COL[2593] = 1'b0;
assign COL[2594] = 1'b0;
assign COL[2595] = 1'b0;
assign COL[2596] = 1'b0;
assign COL[2597] = 1'b0;
assign COL[2598] = 1'b0;
assign COL[2599] = 1'b0;
assign COL[2600] = 1'b1;
assign COL[2601] = 1'b1;
assign COL[2602] = 1'b1;
assign COL[2603] = 1'b1;
assign COL[2604] = 1'b0;
assign COL[2605] = 1'b0;
assign COL[2606] = 1'b0;
assign COL[2607] = 1'b0;
assign COL[2608] = 1'b0;
assign COL[2609] = 1'b0;
assign COL[2610] = 1'b0;
assign COL[2611] = 1'b0;
assign COL[2612] = 1'b0;
assign COL[2613] = 1'b0;
assign COL[2614] = 1'b0;
assign COL[2615] = 1'b0;
assign COL[2616] = 1'b0;
assign COL[2617] = 1'b0;
assign COL[2618] = 1'b0;
assign COL[2619] = 1'b0;
assign COL[2620] = 1'b0;
assign COL[2621] = 1'b0;
assign COL[2622] = 1'b0;
assign COL[2623] = 1'b0;
assign COL[2624] = 1'b0;
assign COL[2625] = 1'b0;
assign COL[2626] = 1'b0;
assign COL[2627] = 1'b0;
assign COL[2628] = 1'b0;
assign COL[2629] = 1'b0;
assign COL[2630] = 1'b0;
assign COL[2631] = 1'b0;
assign COL[2632] = 1'b1;
assign COL[2633] = 1'b1;
assign COL[2634] = 1'b1;
assign COL[2635] = 1'b1;
assign COL[2636] = 1'b0;
assign COL[2637] = 1'b0;
assign COL[2638] = 1'b0;
assign COL[2639] = 1'b0;
assign COL[2640] = 1'b0;
assign COL[2641] = 1'b0;
assign COL[2642] = 1'b0;
assign COL[2643] = 1'b0;
assign COL[2644] = 1'b0;
assign COL[2645] = 1'b0;
assign COL[2646] = 1'b0;
assign COL[2647] = 1'b0;
assign COL[2648] = 1'b0;
assign COL[2649] = 1'b0;
assign COL[2650] = 1'b1;
assign COL[2651] = 1'b1;
assign COL[2652] = 1'b1;
assign COL[2653] = 1'b1;
assign COL[2654] = 1'b1;
assign COL[2655] = 1'b0;
assign COL[2656] = 1'b0;
assign COL[2657] = 1'b0;
assign COL[2658] = 1'b0;
assign COL[2659] = 1'b0;
assign COL[2660] = 1'b0;
assign COL[2661] = 1'b0;
assign COL[2662] = 1'b0;
assign COL[2663] = 1'b0;
assign COL[2664] = 1'b0;
assign COL[2665] = 1'b0;
assign COL[2666] = 1'b0;
assign COL[2667] = 1'b0;
assign COL[2668] = 1'b0;
assign COL[2669] = 1'b0;
assign COL[2670] = 1'b0;
assign COL[2671] = 1'b0;
assign COL[2672] = 1'b0;
assign COL[2673] = 1'b0;
assign COL[2674] = 1'b0;
assign COL[2675] = 1'b0;
assign COL[2676] = 1'b0;
assign COL[2677] = 1'b0;
assign COL[2678] = 1'b0;
assign COL[2679] = 1'b0;
assign COL[2680] = 1'b0;
assign COL[2681] = 1'b0;
assign COL[2682] = 1'b0;
assign COL[2683] = 1'b0;
assign COL[2684] = 1'b0;
assign COL[2685] = 1'b0;
assign COL[2686] = 1'b0;
assign COL[2687] = 1'b0;
assign COL[2688] = 1'b0;
assign COL[2689] = 1'b0;
assign COL[2690] = 1'b0;
assign COL[2691] = 1'b0;
assign COL[2692] = 1'b0;
assign COL[2693] = 1'b0;
assign COL[2694] = 1'b0;
assign COL[2695] = 1'b0;
assign COL[2696] = 1'b0;
assign COL[2697] = 1'b0;
assign COL[2698] = 1'b0;
assign COL[2699] = 1'b0;
assign COL[2700] = 1'b0;
assign COL[2701] = 1'b0;
assign COL[2702] = 1'b0;
assign COL[2703] = 1'b0;
assign COL[2704] = 1'b0;
assign COL[2705] = 1'b0;
assign COL[2706] = 1'b0;
assign COL[2707] = 1'b0;
assign COL[2708] = 1'b0;
assign COL[2709] = 1'b0;
assign COL[2710] = 1'b0;
assign COL[2711] = 1'b0;
assign COL[2712] = 1'b0;
assign COL[2713] = 1'b0;
assign COL[2714] = 1'b0;
assign COL[2715] = 1'b0;
assign COL[2716] = 1'b0;
assign COL[2717] = 1'b0;
assign COL[2718] = 1'b0;
assign COL[2719] = 1'b0;
assign COL[2720] = 1'b0;
assign COL[2721] = 1'b1;
assign COL[2722] = 1'b1;
assign COL[2723] = 1'b1;
assign COL[2724] = 1'b1;
assign COL[2725] = 1'b1;
assign COL[2726] = 1'b0;
assign COL[2727] = 1'b0;
assign COL[2728] = 1'b0;
assign COL[2729] = 1'b0;
assign COL[2730] = 1'b0;
assign COL[2731] = 1'b0;
assign COL[2732] = 1'b0;
assign COL[2733] = 1'b0;
assign COL[2734] = 1'b0;
assign COL[2735] = 1'b0;
assign COL[2736] = 1'b0;
assign COL[2737] = 1'b0;
assign COL[2738] = 1'b0;
assign COL[2739] = 1'b0;
assign COL[2740] = 1'b0;
assign COL[2741] = 1'b0;
assign COL[2742] = 1'b0;
assign COL[2743] = 1'b0;
assign COL[2744] = 1'b0;
assign COL[2745] = 1'b0;
assign COL[2746] = 1'b0;
assign COL[2747] = 1'b0;
assign COL[2748] = 1'b0;
assign COL[2749] = 1'b0;
assign COL[2750] = 1'b0;
assign COL[2751] = 1'b0;
assign COL[2752] = 1'b0;
assign COL[2753] = 1'b0;
assign COL[2754] = 1'b0;
assign COL[2755] = 1'b0;
assign COL[2756] = 1'b0;
assign COL[2757] = 1'b0;
assign COL[2758] = 1'b0;
assign COL[2759] = 1'b0;
assign COL[2760] = 1'b1;
assign COL[2761] = 1'b1;
assign COL[2762] = 1'b1;
assign COL[2763] = 1'b1;
assign COL[2764] = 1'b0;
assign COL[2765] = 1'b0;
assign COL[2766] = 1'b0;
assign COL[2767] = 1'b0;
assign COL[2768] = 1'b0;
assign COL[2769] = 1'b0;
assign COL[2770] = 1'b0;
assign COL[2771] = 1'b0;
assign COL[2772] = 1'b0;
assign COL[2773] = 1'b0;
assign COL[2774] = 1'b0;
assign COL[2775] = 1'b0;
assign COL[2776] = 1'b0;
assign COL[2777] = 1'b0;
assign COL[2778] = 1'b0;
assign COL[2779] = 1'b0;
assign COL[2780] = 1'b0;
assign COL[2781] = 1'b0;
assign COL[2782] = 1'b0;
assign COL[2783] = 1'b0;
assign COL[2784] = 1'b0;
assign COL[2785] = 1'b0;
assign COL[2786] = 1'b0;
assign COL[2787] = 1'b0;
assign COL[2788] = 1'b0;
assign COL[2789] = 1'b0;
assign COL[2790] = 1'b0;
assign COL[2791] = 1'b0;
assign COL[2792] = 1'b1;
assign COL[2793] = 1'b1;
assign COL[2794] = 1'b1;
assign COL[2795] = 1'b1;
assign COL[2796] = 1'b0;
assign COL[2797] = 1'b0;
assign COL[2798] = 1'b0;
assign COL[2799] = 1'b0;
assign COL[2800] = 1'b0;
assign COL[2801] = 1'b0;
assign COL[2802] = 1'b0;
assign COL[2803] = 1'b0;
assign COL[2804] = 1'b0;
assign COL[2805] = 1'b0;
assign COL[2806] = 1'b0;
assign COL[2807] = 1'b0;
assign COL[2808] = 1'b0;
assign COL[2809] = 1'b0;
assign COL[2810] = 1'b1;
assign COL[2811] = 1'b1;
assign COL[2812] = 1'b1;
assign COL[2813] = 1'b1;
assign COL[2814] = 1'b1;
assign COL[2815] = 1'b0;
assign COL[2816] = 1'b0;
assign COL[2817] = 1'b0;
assign COL[2818] = 1'b0;
assign COL[2819] = 1'b0;
assign COL[2820] = 1'b0;
assign COL[2821] = 1'b0;
assign COL[2822] = 1'b0;
assign COL[2823] = 1'b0;
assign COL[2824] = 1'b0;
assign COL[2825] = 1'b0;
assign COL[2826] = 1'b0;
assign COL[2827] = 1'b0;
assign COL[2828] = 1'b0;
assign COL[2829] = 1'b0;
assign COL[2830] = 1'b0;
assign COL[2831] = 1'b0;
assign COL[2832] = 1'b0;
assign COL[2833] = 1'b0;
assign COL[2834] = 1'b0;
assign COL[2835] = 1'b0;
assign COL[2836] = 1'b0;
assign COL[2837] = 1'b0;
assign COL[2838] = 1'b0;
assign COL[2839] = 1'b0;
assign COL[2840] = 1'b0;
assign COL[2841] = 1'b0;
assign COL[2842] = 1'b0;
assign COL[2843] = 1'b0;
assign COL[2844] = 1'b0;
assign COL[2845] = 1'b0;
assign COL[2846] = 1'b0;
assign COL[2847] = 1'b0;
assign COL[2848] = 1'b0;
assign COL[2849] = 1'b0;
assign COL[2850] = 1'b0;
assign COL[2851] = 1'b0;
assign COL[2852] = 1'b0;
assign COL[2853] = 1'b0;
assign COL[2854] = 1'b0;
assign COL[2855] = 1'b0;
assign COL[2856] = 1'b0;
assign COL[2857] = 1'b0;
assign COL[2858] = 1'b0;
assign COL[2859] = 1'b0;
assign COL[2860] = 1'b0;
assign COL[2861] = 1'b0;
assign COL[2862] = 1'b0;
assign COL[2863] = 1'b0;
assign COL[2864] = 1'b0;
assign COL[2865] = 1'b0;
assign COL[2866] = 1'b0;
assign COL[2867] = 1'b0;
assign COL[2868] = 1'b0;
assign COL[2869] = 1'b0;
assign COL[2870] = 1'b0;
assign COL[2871] = 1'b0;
assign COL[2872] = 1'b0;
assign COL[2873] = 1'b0;
assign COL[2874] = 1'b0;
assign COL[2875] = 1'b0;
assign COL[2876] = 1'b0;
assign COL[2877] = 1'b0;
assign COL[2878] = 1'b0;
assign COL[2879] = 1'b0;
assign COL[2880] = 1'b0;
assign COL[2881] = 1'b1;
assign COL[2882] = 1'b1;
assign COL[2883] = 1'b1;
assign COL[2884] = 1'b1;
assign COL[2885] = 1'b1;
assign COL[2886] = 1'b0;
assign COL[2887] = 1'b0;
assign COL[2888] = 1'b0;
assign COL[2889] = 1'b0;
assign COL[2890] = 1'b0;
assign COL[2891] = 1'b0;
assign COL[2892] = 1'b0;
assign COL[2893] = 1'b0;
assign COL[2894] = 1'b0;
assign COL[2895] = 1'b0;
assign COL[2896] = 1'b0;
assign COL[2897] = 1'b0;
assign COL[2898] = 1'b0;
assign COL[2899] = 1'b0;
assign COL[2900] = 1'b0;
assign COL[2901] = 1'b0;
assign COL[2902] = 1'b0;
assign COL[2903] = 1'b0;
assign COL[2904] = 1'b0;
assign COL[2905] = 1'b0;
assign COL[2906] = 1'b0;
assign COL[2907] = 1'b0;
assign COL[2908] = 1'b0;
assign COL[2909] = 1'b0;
assign COL[2910] = 1'b0;
assign COL[2911] = 1'b0;
assign COL[2912] = 1'b0;
assign COL[2913] = 1'b0;
assign COL[2914] = 1'b0;
assign COL[2915] = 1'b0;
assign COL[2916] = 1'b0;
assign COL[2917] = 1'b0;
assign COL[2918] = 1'b0;
assign COL[2919] = 1'b0;
assign COL[2920] = 1'b1;
assign COL[2921] = 1'b1;
assign COL[2922] = 1'b1;
assign COL[2923] = 1'b1;
assign COL[2924] = 1'b0;
assign COL[2925] = 1'b0;
assign COL[2926] = 1'b0;
assign COL[2927] = 1'b0;
assign COL[2928] = 1'b0;
assign COL[2929] = 1'b0;
assign COL[2930] = 1'b0;
assign COL[2931] = 1'b0;
assign COL[2932] = 1'b0;
assign COL[2933] = 1'b0;
assign COL[2934] = 1'b0;
assign COL[2935] = 1'b0;
assign COL[2936] = 1'b0;
assign COL[2937] = 1'b0;
assign COL[2938] = 1'b0;
assign COL[2939] = 1'b0;
assign COL[2940] = 1'b0;
assign COL[2941] = 1'b0;
assign COL[2942] = 1'b0;
assign COL[2943] = 1'b0;
assign COL[2944] = 1'b0;
assign COL[2945] = 1'b0;
assign COL[2946] = 1'b0;
assign COL[2947] = 1'b0;
assign COL[2948] = 1'b0;
assign COL[2949] = 1'b0;
assign COL[2950] = 1'b0;
assign COL[2951] = 1'b0;
assign COL[2952] = 1'b1;
assign COL[2953] = 1'b1;
assign COL[2954] = 1'b1;
assign COL[2955] = 1'b1;
assign COL[2956] = 1'b0;
assign COL[2957] = 1'b0;
assign COL[2958] = 1'b0;
assign COL[2959] = 1'b0;
assign COL[2960] = 1'b0;
assign COL[2961] = 1'b0;
assign COL[2962] = 1'b0;
assign COL[2963] = 1'b0;
assign COL[2964] = 1'b0;
assign COL[2965] = 1'b0;
assign COL[2966] = 1'b0;
assign COL[2967] = 1'b0;
assign COL[2968] = 1'b0;
assign COL[2969] = 1'b0;
assign COL[2970] = 1'b1;
assign COL[2971] = 1'b1;
assign COL[2972] = 1'b1;
assign COL[2973] = 1'b1;
assign COL[2974] = 1'b1;
assign COL[2975] = 1'b0;
assign COL[2976] = 1'b0;
assign COL[2977] = 1'b0;
assign COL[2978] = 1'b0;
assign COL[2979] = 1'b0;
assign COL[2980] = 1'b0;
assign COL[2981] = 1'b0;
assign COL[2982] = 1'b0;
assign COL[2983] = 1'b0;
assign COL[2984] = 1'b0;
assign COL[2985] = 1'b0;
assign COL[2986] = 1'b0;
assign COL[2987] = 1'b0;
assign COL[2988] = 1'b0;
assign COL[2989] = 1'b0;
assign COL[2990] = 1'b0;
assign COL[2991] = 1'b0;
assign COL[2992] = 1'b0;
assign COL[2993] = 1'b0;
assign COL[2994] = 1'b0;
assign COL[2995] = 1'b0;
assign COL[2996] = 1'b0;
assign COL[2997] = 1'b0;
assign COL[2998] = 1'b0;
assign COL[2999] = 1'b0;
assign COL[3000] = 1'b0;
assign COL[3001] = 1'b0;
assign COL[3002] = 1'b0;
assign COL[3003] = 1'b0;
assign COL[3004] = 1'b0;
assign COL[3005] = 1'b0;
assign COL[3006] = 1'b0;
assign COL[3007] = 1'b0;
assign COL[3008] = 1'b0;
assign COL[3009] = 1'b0;
assign COL[3010] = 1'b0;
assign COL[3011] = 1'b0;
assign COL[3012] = 1'b0;
assign COL[3013] = 1'b0;
assign COL[3014] = 1'b0;
assign COL[3015] = 1'b0;
assign COL[3016] = 1'b0;
assign COL[3017] = 1'b0;
assign COL[3018] = 1'b0;
assign COL[3019] = 1'b0;
assign COL[3020] = 1'b0;
assign COL[3021] = 1'b0;
assign COL[3022] = 1'b0;
assign COL[3023] = 1'b0;
assign COL[3024] = 1'b0;
assign COL[3025] = 1'b0;
assign COL[3026] = 1'b0;
assign COL[3027] = 1'b0;
assign COL[3028] = 1'b0;
assign COL[3029] = 1'b0;
assign COL[3030] = 1'b0;
assign COL[3031] = 1'b0;
assign COL[3032] = 1'b0;
assign COL[3033] = 1'b0;
assign COL[3034] = 1'b0;
assign COL[3035] = 1'b0;
assign COL[3036] = 1'b0;
assign COL[3037] = 1'b0;
assign COL[3038] = 1'b0;
assign COL[3039] = 1'b0;
assign COL[3040] = 1'b0;
assign COL[3041] = 1'b1;
assign COL[3042] = 1'b1;
assign COL[3043] = 1'b1;
assign COL[3044] = 1'b1;
assign COL[3045] = 1'b1;
assign COL[3046] = 1'b0;
assign COL[3047] = 1'b0;
assign COL[3048] = 1'b0;
assign COL[3049] = 1'b0;
assign COL[3050] = 1'b0;
assign COL[3051] = 1'b0;
assign COL[3052] = 1'b0;
assign COL[3053] = 1'b0;
assign COL[3054] = 1'b0;
assign COL[3055] = 1'b0;
assign COL[3056] = 1'b0;
assign COL[3057] = 1'b0;
assign COL[3058] = 1'b0;
assign COL[3059] = 1'b0;
assign COL[3060] = 1'b0;
assign COL[3061] = 1'b0;
assign COL[3062] = 1'b0;
assign COL[3063] = 1'b0;
assign COL[3064] = 1'b0;
assign COL[3065] = 1'b0;
assign COL[3066] = 1'b0;
assign COL[3067] = 1'b0;
assign COL[3068] = 1'b0;
assign COL[3069] = 1'b0;
assign COL[3070] = 1'b0;
assign COL[3071] = 1'b0;
assign COL[3072] = 1'b0;
assign COL[3073] = 1'b0;
assign COL[3074] = 1'b0;
assign COL[3075] = 1'b0;
assign COL[3076] = 1'b0;
assign COL[3077] = 1'b0;
assign COL[3078] = 1'b0;
assign COL[3079] = 1'b0;
assign COL[3080] = 1'b1;
assign COL[3081] = 1'b1;
assign COL[3082] = 1'b1;
assign COL[3083] = 1'b1;
assign COL[3084] = 1'b0;
assign COL[3085] = 1'b0;
assign COL[3086] = 1'b0;
assign COL[3087] = 1'b0;
assign COL[3088] = 1'b0;
assign COL[3089] = 1'b0;
assign COL[3090] = 1'b0;
assign COL[3091] = 1'b0;
assign COL[3092] = 1'b0;
assign COL[3093] = 1'b0;
assign COL[3094] = 1'b0;
assign COL[3095] = 1'b0;
assign COL[3096] = 1'b0;
assign COL[3097] = 1'b0;
assign COL[3098] = 1'b0;
assign COL[3099] = 1'b0;
assign COL[3100] = 1'b0;
assign COL[3101] = 1'b0;
assign COL[3102] = 1'b0;
assign COL[3103] = 1'b0;
assign COL[3104] = 1'b0;
assign COL[3105] = 1'b0;
assign COL[3106] = 1'b0;
assign COL[3107] = 1'b0;
assign COL[3108] = 1'b0;
assign COL[3109] = 1'b0;
assign COL[3110] = 1'b0;
assign COL[3111] = 1'b0;
assign COL[3112] = 1'b1;
assign COL[3113] = 1'b1;
assign COL[3114] = 1'b1;
assign COL[3115] = 1'b1;
assign COL[3116] = 1'b0;
assign COL[3117] = 1'b0;
assign COL[3118] = 1'b0;
assign COL[3119] = 1'b0;
assign COL[3120] = 1'b0;
assign COL[3121] = 1'b0;
assign COL[3122] = 1'b0;
assign COL[3123] = 1'b0;
assign COL[3124] = 1'b0;
assign COL[3125] = 1'b0;
assign COL[3126] = 1'b0;
assign COL[3127] = 1'b0;
assign COL[3128] = 1'b0;
assign COL[3129] = 1'b0;
assign COL[3130] = 1'b1;
assign COL[3131] = 1'b1;
assign COL[3132] = 1'b1;
assign COL[3133] = 1'b1;
assign COL[3134] = 1'b1;
assign COL[3135] = 1'b0;
assign COL[3136] = 1'b0;
assign COL[3137] = 1'b0;
assign COL[3138] = 1'b0;
assign COL[3139] = 1'b0;
assign COL[3140] = 1'b0;
assign COL[3141] = 1'b0;
assign COL[3142] = 1'b0;
assign COL[3143] = 1'b0;
assign COL[3144] = 1'b0;
assign COL[3145] = 1'b0;
assign COL[3146] = 1'b0;
assign COL[3147] = 1'b0;
assign COL[3148] = 1'b0;
assign COL[3149] = 1'b0;
assign COL[3150] = 1'b0;
assign COL[3151] = 1'b0;
assign COL[3152] = 1'b0;
assign COL[3153] = 1'b0;
assign COL[3154] = 1'b0;
assign COL[3155] = 1'b0;
assign COL[3156] = 1'b0;
assign COL[3157] = 1'b0;
assign COL[3158] = 1'b0;
assign COL[3159] = 1'b0;
assign COL[3160] = 1'b0;
assign COL[3161] = 1'b0;
assign COL[3162] = 1'b0;
assign COL[3163] = 1'b0;
assign COL[3164] = 1'b0;
assign COL[3165] = 1'b0;
assign COL[3166] = 1'b0;
assign COL[3167] = 1'b0;
assign COL[3168] = 1'b0;
assign COL[3169] = 1'b0;
assign COL[3170] = 1'b0;
assign COL[3171] = 1'b0;
assign COL[3172] = 1'b0;
assign COL[3173] = 1'b0;
assign COL[3174] = 1'b0;
assign COL[3175] = 1'b0;
assign COL[3176] = 1'b0;
assign COL[3177] = 1'b0;
assign COL[3178] = 1'b0;
assign COL[3179] = 1'b0;
assign COL[3180] = 1'b0;
assign COL[3181] = 1'b0;
assign COL[3182] = 1'b0;
assign COL[3183] = 1'b0;
assign COL[3184] = 1'b0;
assign COL[3185] = 1'b0;
assign COL[3186] = 1'b0;
assign COL[3187] = 1'b0;
assign COL[3188] = 1'b0;
assign COL[3189] = 1'b0;
assign COL[3190] = 1'b0;
assign COL[3191] = 1'b0;
assign COL[3192] = 1'b0;
assign COL[3193] = 1'b0;
assign COL[3194] = 1'b0;
assign COL[3195] = 1'b0;
assign COL[3196] = 1'b0;
assign COL[3197] = 1'b0;
assign COL[3198] = 1'b0;
assign COL[3199] = 1'b0;
assign COL[3200] = 1'b0;
assign COL[3201] = 1'b1;
assign COL[3202] = 1'b1;
assign COL[3203] = 1'b1;
assign COL[3204] = 1'b1;
assign COL[3205] = 1'b1;
assign COL[3206] = 1'b0;
assign COL[3207] = 1'b0;
assign COL[3208] = 1'b0;
assign COL[3209] = 1'b0;
assign COL[3210] = 1'b0;
assign COL[3211] = 1'b0;
assign COL[3212] = 1'b0;
assign COL[3213] = 1'b0;
assign COL[3214] = 1'b0;
assign COL[3215] = 1'b0;
assign COL[3216] = 1'b1;
assign COL[3217] = 1'b1;
assign COL[3218] = 1'b1;
assign COL[3219] = 1'b1;
assign COL[3220] = 1'b1;
assign COL[3221] = 1'b1;
assign COL[3222] = 1'b1;
assign COL[3223] = 1'b1;
assign COL[3224] = 1'b1;
assign COL[3225] = 1'b1;
assign COL[3226] = 1'b1;
assign COL[3227] = 1'b1;
assign COL[3228] = 1'b1;
assign COL[3229] = 1'b1;
assign COL[3230] = 1'b1;
assign COL[3231] = 1'b1;
assign COL[3232] = 1'b0;
assign COL[3233] = 1'b0;
assign COL[3234] = 1'b0;
assign COL[3235] = 1'b0;
assign COL[3236] = 1'b0;
assign COL[3237] = 1'b0;
assign COL[3238] = 1'b0;
assign COL[3239] = 1'b0;
assign COL[3240] = 1'b1;
assign COL[3241] = 1'b1;
assign COL[3242] = 1'b1;
assign COL[3243] = 1'b1;
assign COL[3244] = 1'b0;
assign COL[3245] = 1'b0;
assign COL[3246] = 1'b0;
assign COL[3247] = 1'b0;
assign COL[3248] = 1'b0;
assign COL[3249] = 1'b0;
assign COL[3250] = 1'b0;
assign COL[3251] = 1'b0;
assign COL[3252] = 1'b0;
assign COL[3253] = 1'b0;
assign COL[3254] = 1'b0;
assign COL[3255] = 1'b0;
assign COL[3256] = 1'b0;
assign COL[3257] = 1'b0;
assign COL[3258] = 1'b0;
assign COL[3259] = 1'b0;
assign COL[3260] = 1'b0;
assign COL[3261] = 1'b0;
assign COL[3262] = 1'b0;
assign COL[3263] = 1'b0;
assign COL[3264] = 1'b0;
assign COL[3265] = 1'b0;
assign COL[3266] = 1'b0;
assign COL[3267] = 1'b0;
assign COL[3268] = 1'b0;
assign COL[3269] = 1'b0;
assign COL[3270] = 1'b0;
assign COL[3271] = 1'b0;
assign COL[3272] = 1'b1;
assign COL[3273] = 1'b1;
assign COL[3274] = 1'b1;
assign COL[3275] = 1'b1;
assign COL[3276] = 1'b0;
assign COL[3277] = 1'b0;
assign COL[3278] = 1'b0;
assign COL[3279] = 1'b0;
assign COL[3280] = 1'b0;
assign COL[3281] = 1'b0;
assign COL[3282] = 1'b0;
assign COL[3283] = 1'b0;
assign COL[3284] = 1'b0;
assign COL[3285] = 1'b0;
assign COL[3286] = 1'b0;
assign COL[3287] = 1'b0;
assign COL[3288] = 1'b0;
assign COL[3289] = 1'b0;
assign COL[3290] = 1'b1;
assign COL[3291] = 1'b1;
assign COL[3292] = 1'b1;
assign COL[3293] = 1'b1;
assign COL[3294] = 1'b1;
assign COL[3295] = 1'b0;
assign COL[3296] = 1'b0;
assign COL[3297] = 1'b0;
assign COL[3298] = 1'b0;
assign COL[3299] = 1'b0;
assign COL[3300] = 1'b0;
assign COL[3301] = 1'b0;
assign COL[3302] = 1'b0;
assign COL[3303] = 1'b0;
assign COL[3304] = 1'b0;
assign COL[3305] = 1'b0;
assign COL[3306] = 1'b0;
assign COL[3307] = 1'b0;
assign COL[3308] = 1'b0;
assign COL[3309] = 1'b0;
assign COL[3310] = 1'b0;
assign COL[3311] = 1'b0;
assign COL[3312] = 1'b0;
assign COL[3313] = 1'b0;
assign COL[3314] = 1'b0;
assign COL[3315] = 1'b0;
assign COL[3316] = 1'b0;
assign COL[3317] = 1'b0;
assign COL[3318] = 1'b0;
assign COL[3319] = 1'b0;
assign COL[3320] = 1'b0;
assign COL[3321] = 1'b0;
assign COL[3322] = 1'b0;
assign COL[3323] = 1'b0;
assign COL[3324] = 1'b0;
assign COL[3325] = 1'b0;
assign COL[3326] = 1'b0;
assign COL[3327] = 1'b0;
assign COL[3328] = 1'b0;
assign COL[3329] = 1'b0;
assign COL[3330] = 1'b0;
assign COL[3331] = 1'b0;
assign COL[3332] = 1'b0;
assign COL[3333] = 1'b0;
assign COL[3334] = 1'b0;
assign COL[3335] = 1'b0;
assign COL[3336] = 1'b0;
assign COL[3337] = 1'b0;
assign COL[3338] = 1'b0;
assign COL[3339] = 1'b0;
assign COL[3340] = 1'b0;
assign COL[3341] = 1'b0;
assign COL[3342] = 1'b0;
assign COL[3343] = 1'b0;
assign COL[3344] = 1'b0;
assign COL[3345] = 1'b0;
assign COL[3346] = 1'b0;
assign COL[3347] = 1'b0;
assign COL[3348] = 1'b0;
assign COL[3349] = 1'b0;
assign COL[3350] = 1'b0;
assign COL[3351] = 1'b0;
assign COL[3352] = 1'b0;
assign COL[3353] = 1'b0;
assign COL[3354] = 1'b0;
assign COL[3355] = 1'b0;
assign COL[3356] = 1'b0;
assign COL[3357] = 1'b0;
assign COL[3358] = 1'b0;
assign COL[3359] = 1'b0;
assign COL[3360] = 1'b0;
assign COL[3361] = 1'b1;
assign COL[3362] = 1'b1;
assign COL[3363] = 1'b1;
assign COL[3364] = 1'b1;
assign COL[3365] = 1'b1;
assign COL[3366] = 1'b0;
assign COL[3367] = 1'b0;
assign COL[3368] = 1'b0;
assign COL[3369] = 1'b0;
assign COL[3370] = 1'b0;
assign COL[3371] = 1'b0;
assign COL[3372] = 1'b0;
assign COL[3373] = 1'b0;
assign COL[3374] = 1'b0;
assign COL[3375] = 1'b0;
assign COL[3376] = 1'b1;
assign COL[3377] = 1'b1;
assign COL[3378] = 1'b1;
assign COL[3379] = 1'b1;
assign COL[3380] = 1'b1;
assign COL[3381] = 1'b1;
assign COL[3382] = 1'b1;
assign COL[3383] = 1'b1;
assign COL[3384] = 1'b1;
assign COL[3385] = 1'b1;
assign COL[3386] = 1'b1;
assign COL[3387] = 1'b1;
assign COL[3388] = 1'b1;
assign COL[3389] = 1'b1;
assign COL[3390] = 1'b1;
assign COL[3391] = 1'b1;
assign COL[3392] = 1'b0;
assign COL[3393] = 1'b0;
assign COL[3394] = 1'b0;
assign COL[3395] = 1'b0;
assign COL[3396] = 1'b0;
assign COL[3397] = 1'b0;
assign COL[3398] = 1'b0;
assign COL[3399] = 1'b0;
assign COL[3400] = 1'b1;
assign COL[3401] = 1'b1;
assign COL[3402] = 1'b1;
assign COL[3403] = 1'b1;
assign COL[3404] = 1'b0;
assign COL[3405] = 1'b0;
assign COL[3406] = 1'b0;
assign COL[3407] = 1'b0;
assign COL[3408] = 1'b0;
assign COL[3409] = 1'b0;
assign COL[3410] = 1'b1;
assign COL[3411] = 1'b1;
assign COL[3412] = 1'b1;
assign COL[3413] = 1'b1;
assign COL[3414] = 1'b1;
assign COL[3415] = 1'b1;
assign COL[3416] = 1'b1;
assign COL[3417] = 1'b1;
assign COL[3418] = 1'b1;
assign COL[3419] = 1'b1;
assign COL[3420] = 1'b1;
assign COL[3421] = 1'b1;
assign COL[3422] = 1'b1;
assign COL[3423] = 1'b1;
assign COL[3424] = 1'b1;
assign COL[3425] = 1'b1;
assign COL[3426] = 1'b0;
assign COL[3427] = 1'b0;
assign COL[3428] = 1'b0;
assign COL[3429] = 1'b0;
assign COL[3430] = 1'b0;
assign COL[3431] = 1'b0;
assign COL[3432] = 1'b1;
assign COL[3433] = 1'b1;
assign COL[3434] = 1'b1;
assign COL[3435] = 1'b1;
assign COL[3436] = 1'b0;
assign COL[3437] = 1'b0;
assign COL[3438] = 1'b0;
assign COL[3439] = 1'b0;
assign COL[3440] = 1'b0;
assign COL[3441] = 1'b0;
assign COL[3442] = 1'b0;
assign COL[3443] = 1'b0;
assign COL[3444] = 1'b0;
assign COL[3445] = 1'b0;
assign COL[3446] = 1'b0;
assign COL[3447] = 1'b0;
assign COL[3448] = 1'b0;
assign COL[3449] = 1'b0;
assign COL[3450] = 1'b1;
assign COL[3451] = 1'b1;
assign COL[3452] = 1'b1;
assign COL[3453] = 1'b1;
assign COL[3454] = 1'b1;
assign COL[3455] = 1'b0;
assign COL[3456] = 1'b0;
assign COL[3457] = 1'b0;
assign COL[3458] = 1'b0;
assign COL[3459] = 1'b0;
assign COL[3460] = 1'b0;
assign COL[3461] = 1'b0;
assign COL[3462] = 1'b0;
assign COL[3463] = 1'b0;
assign COL[3464] = 1'b0;
assign COL[3465] = 1'b0;
assign COL[3466] = 1'b0;
assign COL[3467] = 1'b0;
assign COL[3468] = 1'b0;
assign COL[3469] = 1'b0;
assign COL[3470] = 1'b0;
assign COL[3471] = 1'b0;
assign COL[3472] = 1'b0;
assign COL[3473] = 1'b0;
assign COL[3474] = 1'b0;
assign COL[3475] = 1'b0;
assign COL[3476] = 1'b0;
assign COL[3477] = 1'b0;
assign COL[3478] = 1'b0;
assign COL[3479] = 1'b0;
assign COL[3480] = 1'b0;
assign COL[3481] = 1'b0;
assign COL[3482] = 1'b0;
assign COL[3483] = 1'b0;
assign COL[3484] = 1'b0;
assign COL[3485] = 1'b0;
assign COL[3486] = 1'b0;
assign COL[3487] = 1'b0;
assign COL[3488] = 1'b0;
assign COL[3489] = 1'b0;
assign COL[3490] = 1'b0;
assign COL[3491] = 1'b0;
assign COL[3492] = 1'b0;
assign COL[3493] = 1'b0;
assign COL[3494] = 1'b0;
assign COL[3495] = 1'b0;
assign COL[3496] = 1'b0;
assign COL[3497] = 1'b0;
assign COL[3498] = 1'b0;
assign COL[3499] = 1'b0;
assign COL[3500] = 1'b0;
assign COL[3501] = 1'b0;
assign COL[3502] = 1'b0;
assign COL[3503] = 1'b0;
assign COL[3504] = 1'b0;
assign COL[3505] = 1'b0;
assign COL[3506] = 1'b0;
assign COL[3507] = 1'b0;
assign COL[3508] = 1'b0;
assign COL[3509] = 1'b0;
assign COL[3510] = 1'b0;
assign COL[3511] = 1'b0;
assign COL[3512] = 1'b0;
assign COL[3513] = 1'b0;
assign COL[3514] = 1'b0;
assign COL[3515] = 1'b0;
assign COL[3516] = 1'b0;
assign COL[3517] = 1'b0;
assign COL[3518] = 1'b0;
assign COL[3519] = 1'b0;
assign COL[3520] = 1'b0;
assign COL[3521] = 1'b1;
assign COL[3522] = 1'b1;
assign COL[3523] = 1'b1;
assign COL[3524] = 1'b1;
assign COL[3525] = 1'b1;
assign COL[3526] = 1'b0;
assign COL[3527] = 1'b0;
assign COL[3528] = 1'b0;
assign COL[3529] = 1'b0;
assign COL[3530] = 1'b0;
assign COL[3531] = 1'b0;
assign COL[3532] = 1'b0;
assign COL[3533] = 1'b0;
assign COL[3534] = 1'b0;
assign COL[3535] = 1'b0;
assign COL[3536] = 1'b1;
assign COL[3537] = 1'b1;
assign COL[3538] = 1'b1;
assign COL[3539] = 1'b1;
assign COL[3540] = 1'b1;
assign COL[3541] = 1'b1;
assign COL[3542] = 1'b1;
assign COL[3543] = 1'b1;
assign COL[3544] = 1'b1;
assign COL[3545] = 1'b1;
assign COL[3546] = 1'b1;
assign COL[3547] = 1'b1;
assign COL[3548] = 1'b1;
assign COL[3549] = 1'b1;
assign COL[3550] = 1'b1;
assign COL[3551] = 1'b1;
assign COL[3552] = 1'b0;
assign COL[3553] = 1'b0;
assign COL[3554] = 1'b0;
assign COL[3555] = 1'b0;
assign COL[3556] = 1'b0;
assign COL[3557] = 1'b0;
assign COL[3558] = 1'b0;
assign COL[3559] = 1'b0;
assign COL[3560] = 1'b1;
assign COL[3561] = 1'b1;
assign COL[3562] = 1'b1;
assign COL[3563] = 1'b1;
assign COL[3564] = 1'b0;
assign COL[3565] = 1'b0;
assign COL[3566] = 1'b0;
assign COL[3567] = 1'b0;
assign COL[3568] = 1'b0;
assign COL[3569] = 1'b0;
assign COL[3570] = 1'b1;
assign COL[3571] = 1'b1;
assign COL[3572] = 1'b1;
assign COL[3573] = 1'b1;
assign COL[3574] = 1'b1;
assign COL[3575] = 1'b1;
assign COL[3576] = 1'b1;
assign COL[3577] = 1'b1;
assign COL[3578] = 1'b1;
assign COL[3579] = 1'b1;
assign COL[3580] = 1'b1;
assign COL[3581] = 1'b1;
assign COL[3582] = 1'b1;
assign COL[3583] = 1'b1;
assign COL[3584] = 1'b1;
assign COL[3585] = 1'b1;
assign COL[3586] = 1'b0;
assign COL[3587] = 1'b0;
assign COL[3588] = 1'b0;
assign COL[3589] = 1'b0;
assign COL[3590] = 1'b0;
assign COL[3591] = 1'b0;
assign COL[3592] = 1'b1;
assign COL[3593] = 1'b1;
assign COL[3594] = 1'b1;
assign COL[3595] = 1'b1;
assign COL[3596] = 1'b0;
assign COL[3597] = 1'b0;
assign COL[3598] = 1'b0;
assign COL[3599] = 1'b0;
assign COL[3600] = 1'b0;
assign COL[3601] = 1'b0;
assign COL[3602] = 1'b0;
assign COL[3603] = 1'b0;
assign COL[3604] = 1'b0;
assign COL[3605] = 1'b0;
assign COL[3606] = 1'b0;
assign COL[3607] = 1'b0;
assign COL[3608] = 1'b0;
assign COL[3609] = 1'b0;
assign COL[3610] = 1'b1;
assign COL[3611] = 1'b1;
assign COL[3612] = 1'b1;
assign COL[3613] = 1'b1;
assign COL[3614] = 1'b1;
assign COL[3615] = 1'b0;
assign COL[3616] = 1'b0;
assign COL[3617] = 1'b0;
assign COL[3618] = 1'b0;
assign COL[3619] = 1'b0;
assign COL[3620] = 1'b0;
assign COL[3621] = 1'b0;
assign COL[3622] = 1'b0;
assign COL[3623] = 1'b0;
assign COL[3624] = 1'b0;
assign COL[3625] = 1'b0;
assign COL[3626] = 1'b0;
assign COL[3627] = 1'b0;
assign COL[3628] = 1'b0;
assign COL[3629] = 1'b0;
assign COL[3630] = 1'b0;
assign COL[3631] = 1'b0;
assign COL[3632] = 1'b0;
assign COL[3633] = 1'b0;
assign COL[3634] = 1'b0;
assign COL[3635] = 1'b0;
assign COL[3636] = 1'b0;
assign COL[3637] = 1'b0;
assign COL[3638] = 1'b0;
assign COL[3639] = 1'b0;
assign COL[3640] = 1'b0;
assign COL[3641] = 1'b0;
assign COL[3642] = 1'b0;
assign COL[3643] = 1'b0;
assign COL[3644] = 1'b0;
assign COL[3645] = 1'b0;
assign COL[3646] = 1'b0;
assign COL[3647] = 1'b0;
assign COL[3648] = 1'b0;
assign COL[3649] = 1'b0;
assign COL[3650] = 1'b0;
assign COL[3651] = 1'b0;
assign COL[3652] = 1'b0;
assign COL[3653] = 1'b0;
assign COL[3654] = 1'b0;
assign COL[3655] = 1'b0;
assign COL[3656] = 1'b0;
assign COL[3657] = 1'b0;
assign COL[3658] = 1'b0;
assign COL[3659] = 1'b0;
assign COL[3660] = 1'b0;
assign COL[3661] = 1'b0;
assign COL[3662] = 1'b0;
assign COL[3663] = 1'b0;
assign COL[3664] = 1'b0;
assign COL[3665] = 1'b0;
assign COL[3666] = 1'b0;
assign COL[3667] = 1'b0;
assign COL[3668] = 1'b0;
assign COL[3669] = 1'b0;
assign COL[3670] = 1'b0;
assign COL[3671] = 1'b0;
assign COL[3672] = 1'b0;
assign COL[3673] = 1'b0;
assign COL[3674] = 1'b0;
assign COL[3675] = 1'b0;
assign COL[3676] = 1'b0;
assign COL[3677] = 1'b0;
assign COL[3678] = 1'b0;
assign COL[3679] = 1'b0;
assign COL[3680] = 1'b0;
assign COL[3681] = 1'b1;
assign COL[3682] = 1'b1;
assign COL[3683] = 1'b1;
assign COL[3684] = 1'b1;
assign COL[3685] = 1'b1;
assign COL[3686] = 1'b0;
assign COL[3687] = 1'b0;
assign COL[3688] = 1'b0;
assign COL[3689] = 1'b0;
assign COL[3690] = 1'b0;
assign COL[3691] = 1'b0;
assign COL[3692] = 1'b0;
assign COL[3693] = 1'b0;
assign COL[3694] = 1'b0;
assign COL[3695] = 1'b0;
assign COL[3696] = 1'b1;
assign COL[3697] = 1'b1;
assign COL[3698] = 1'b1;
assign COL[3699] = 1'b1;
assign COL[3700] = 1'b1;
assign COL[3701] = 1'b1;
assign COL[3702] = 1'b1;
assign COL[3703] = 1'b1;
assign COL[3704] = 1'b1;
assign COL[3705] = 1'b1;
assign COL[3706] = 1'b1;
assign COL[3707] = 1'b1;
assign COL[3708] = 1'b1;
assign COL[3709] = 1'b1;
assign COL[3710] = 1'b1;
assign COL[3711] = 1'b1;
assign COL[3712] = 1'b0;
assign COL[3713] = 1'b0;
assign COL[3714] = 1'b0;
assign COL[3715] = 1'b0;
assign COL[3716] = 1'b0;
assign COL[3717] = 1'b0;
assign COL[3718] = 1'b0;
assign COL[3719] = 1'b0;
assign COL[3720] = 1'b1;
assign COL[3721] = 1'b1;
assign COL[3722] = 1'b1;
assign COL[3723] = 1'b1;
assign COL[3724] = 1'b0;
assign COL[3725] = 1'b0;
assign COL[3726] = 1'b0;
assign COL[3727] = 1'b0;
assign COL[3728] = 1'b0;
assign COL[3729] = 1'b0;
assign COL[3730] = 1'b1;
assign COL[3731] = 1'b1;
assign COL[3732] = 1'b1;
assign COL[3733] = 1'b1;
assign COL[3734] = 1'b1;
assign COL[3735] = 1'b1;
assign COL[3736] = 1'b1;
assign COL[3737] = 1'b1;
assign COL[3738] = 1'b1;
assign COL[3739] = 1'b1;
assign COL[3740] = 1'b1;
assign COL[3741] = 1'b1;
assign COL[3742] = 1'b1;
assign COL[3743] = 1'b1;
assign COL[3744] = 1'b1;
assign COL[3745] = 1'b1;
assign COL[3746] = 1'b0;
assign COL[3747] = 1'b0;
assign COL[3748] = 1'b0;
assign COL[3749] = 1'b0;
assign COL[3750] = 1'b0;
assign COL[3751] = 1'b0;
assign COL[3752] = 1'b0;
assign COL[3753] = 1'b0;
assign COL[3754] = 1'b0;
assign COL[3755] = 1'b0;
assign COL[3756] = 1'b0;
assign COL[3757] = 1'b0;
assign COL[3758] = 1'b0;
assign COL[3759] = 1'b0;
assign COL[3760] = 1'b0;
assign COL[3761] = 1'b0;
assign COL[3762] = 1'b0;
assign COL[3763] = 1'b0;
assign COL[3764] = 1'b0;
assign COL[3765] = 1'b0;
assign COL[3766] = 1'b0;
assign COL[3767] = 1'b0;
assign COL[3768] = 1'b0;
assign COL[3769] = 1'b0;
assign COL[3770] = 1'b1;
assign COL[3771] = 1'b1;
assign COL[3772] = 1'b1;
assign COL[3773] = 1'b1;
assign COL[3774] = 1'b1;
assign COL[3775] = 1'b0;
assign COL[3776] = 1'b0;
assign COL[3777] = 1'b0;
assign COL[3778] = 1'b0;
assign COL[3779] = 1'b0;
assign COL[3780] = 1'b0;
assign COL[3781] = 1'b0;
assign COL[3782] = 1'b0;
assign COL[3783] = 1'b0;
assign COL[3784] = 1'b0;
assign COL[3785] = 1'b0;
assign COL[3786] = 1'b0;
assign COL[3787] = 1'b0;
assign COL[3788] = 1'b0;
assign COL[3789] = 1'b0;
assign COL[3790] = 1'b0;
assign COL[3791] = 1'b0;
assign COL[3792] = 1'b0;
assign COL[3793] = 1'b0;
assign COL[3794] = 1'b0;
assign COL[3795] = 1'b0;
assign COL[3796] = 1'b0;
assign COL[3797] = 1'b0;
assign COL[3798] = 1'b0;
assign COL[3799] = 1'b0;
assign COL[3800] = 1'b0;
assign COL[3801] = 1'b0;
assign COL[3802] = 1'b0;
assign COL[3803] = 1'b0;
assign COL[3804] = 1'b0;
assign COL[3805] = 1'b0;
assign COL[3806] = 1'b0;
assign COL[3807] = 1'b0;
assign COL[3808] = 1'b0;
assign COL[3809] = 1'b0;
assign COL[3810] = 1'b0;
assign COL[3811] = 1'b0;
assign COL[3812] = 1'b0;
assign COL[3813] = 1'b0;
assign COL[3814] = 1'b0;
assign COL[3815] = 1'b0;
assign COL[3816] = 1'b0;
assign COL[3817] = 1'b0;
assign COL[3818] = 1'b0;
assign COL[3819] = 1'b0;
assign COL[3820] = 1'b0;
assign COL[3821] = 1'b0;
assign COL[3822] = 1'b0;
assign COL[3823] = 1'b0;
assign COL[3824] = 1'b0;
assign COL[3825] = 1'b0;
assign COL[3826] = 1'b0;
assign COL[3827] = 1'b0;
assign COL[3828] = 1'b0;
assign COL[3829] = 1'b0;
assign COL[3830] = 1'b0;
assign COL[3831] = 1'b0;
assign COL[3832] = 1'b0;
assign COL[3833] = 1'b0;
assign COL[3834] = 1'b0;
assign COL[3835] = 1'b0;
assign COL[3836] = 1'b0;
assign COL[3837] = 1'b0;
assign COL[3838] = 1'b0;
assign COL[3839] = 1'b0;
assign COL[3840] = 1'b0;
assign COL[3841] = 1'b1;
assign COL[3842] = 1'b1;
assign COL[3843] = 1'b1;
assign COL[3844] = 1'b1;
assign COL[3845] = 1'b1;
assign COL[3846] = 1'b0;
assign COL[3847] = 1'b0;
assign COL[3848] = 1'b0;
assign COL[3849] = 1'b0;
assign COL[3850] = 1'b0;
assign COL[3851] = 1'b0;
assign COL[3852] = 1'b0;
assign COL[3853] = 1'b0;
assign COL[3854] = 1'b0;
assign COL[3855] = 1'b0;
assign COL[3856] = 1'b1;
assign COL[3857] = 1'b1;
assign COL[3858] = 1'b1;
assign COL[3859] = 1'b1;
assign COL[3860] = 1'b1;
assign COL[3861] = 1'b1;
assign COL[3862] = 1'b1;
assign COL[3863] = 1'b1;
assign COL[3864] = 1'b1;
assign COL[3865] = 1'b1;
assign COL[3866] = 1'b1;
assign COL[3867] = 1'b1;
assign COL[3868] = 1'b1;
assign COL[3869] = 1'b1;
assign COL[3870] = 1'b1;
assign COL[3871] = 1'b1;
assign COL[3872] = 1'b0;
assign COL[3873] = 1'b0;
assign COL[3874] = 1'b0;
assign COL[3875] = 1'b0;
assign COL[3876] = 1'b0;
assign COL[3877] = 1'b0;
assign COL[3878] = 1'b0;
assign COL[3879] = 1'b0;
assign COL[3880] = 1'b1;
assign COL[3881] = 1'b1;
assign COL[3882] = 1'b1;
assign COL[3883] = 1'b1;
assign COL[3884] = 1'b0;
assign COL[3885] = 1'b0;
assign COL[3886] = 1'b0;
assign COL[3887] = 1'b0;
assign COL[3888] = 1'b0;
assign COL[3889] = 1'b0;
assign COL[3890] = 1'b1;
assign COL[3891] = 1'b1;
assign COL[3892] = 1'b1;
assign COL[3893] = 1'b1;
assign COL[3894] = 1'b1;
assign COL[3895] = 1'b1;
assign COL[3896] = 1'b1;
assign COL[3897] = 1'b1;
assign COL[3898] = 1'b1;
assign COL[3899] = 1'b1;
assign COL[3900] = 1'b1;
assign COL[3901] = 1'b1;
assign COL[3902] = 1'b1;
assign COL[3903] = 1'b1;
assign COL[3904] = 1'b1;
assign COL[3905] = 1'b1;
assign COL[3906] = 1'b0;
assign COL[3907] = 1'b0;
assign COL[3908] = 1'b0;
assign COL[3909] = 1'b0;
assign COL[3910] = 1'b0;
assign COL[3911] = 1'b0;
assign COL[3912] = 1'b0;
assign COL[3913] = 1'b0;
assign COL[3914] = 1'b0;
assign COL[3915] = 1'b0;
assign COL[3916] = 1'b0;
assign COL[3917] = 1'b0;
assign COL[3918] = 1'b0;
assign COL[3919] = 1'b0;
assign COL[3920] = 1'b0;
assign COL[3921] = 1'b0;
assign COL[3922] = 1'b0;
assign COL[3923] = 1'b0;
assign COL[3924] = 1'b0;
assign COL[3925] = 1'b0;
assign COL[3926] = 1'b0;
assign COL[3927] = 1'b0;
assign COL[3928] = 1'b0;
assign COL[3929] = 1'b0;
assign COL[3930] = 1'b1;
assign COL[3931] = 1'b1;
assign COL[3932] = 1'b1;
assign COL[3933] = 1'b1;
assign COL[3934] = 1'b1;
assign COL[3935] = 1'b0;
assign COL[3936] = 1'b0;
assign COL[3937] = 1'b0;
assign COL[3938] = 1'b0;
assign COL[3939] = 1'b0;
assign COL[3940] = 1'b0;
assign COL[3941] = 1'b0;
assign COL[3942] = 1'b0;
assign COL[3943] = 1'b0;
assign COL[3944] = 1'b0;
assign COL[3945] = 1'b0;
assign COL[3946] = 1'b0;
assign COL[3947] = 1'b0;
assign COL[3948] = 1'b0;
assign COL[3949] = 1'b0;
assign COL[3950] = 1'b0;
assign COL[3951] = 1'b0;
assign COL[3952] = 1'b0;
assign COL[3953] = 1'b0;
assign COL[3954] = 1'b0;
assign COL[3955] = 1'b0;
assign COL[3956] = 1'b0;
assign COL[3957] = 1'b0;
assign COL[3958] = 1'b0;
assign COL[3959] = 1'b0;
assign COL[3960] = 1'b0;
assign COL[3961] = 1'b0;
assign COL[3962] = 1'b0;
assign COL[3963] = 1'b0;
assign COL[3964] = 1'b0;
assign COL[3965] = 1'b0;
assign COL[3966] = 1'b0;
assign COL[3967] = 1'b0;
assign COL[3968] = 1'b0;
assign COL[3969] = 1'b0;
assign COL[3970] = 1'b0;
assign COL[3971] = 1'b0;
assign COL[3972] = 1'b0;
assign COL[3973] = 1'b0;
assign COL[3974] = 1'b0;
assign COL[3975] = 1'b0;
assign COL[3976] = 1'b0;
assign COL[3977] = 1'b0;
assign COL[3978] = 1'b0;
assign COL[3979] = 1'b0;
assign COL[3980] = 1'b0;
assign COL[3981] = 1'b0;
assign COL[3982] = 1'b0;
assign COL[3983] = 1'b0;
assign COL[3984] = 1'b0;
assign COL[3985] = 1'b0;
assign COL[3986] = 1'b0;
assign COL[3987] = 1'b0;
assign COL[3988] = 1'b0;
assign COL[3989] = 1'b0;
assign COL[3990] = 1'b0;
assign COL[3991] = 1'b0;
assign COL[3992] = 1'b0;
assign COL[3993] = 1'b0;
assign COL[3994] = 1'b0;
assign COL[3995] = 1'b0;
assign COL[3996] = 1'b0;
assign COL[3997] = 1'b0;
assign COL[3998] = 1'b0;
assign COL[3999] = 1'b0;
assign COL[4000] = 1'b0;
assign COL[4001] = 1'b1;
assign COL[4002] = 1'b1;
assign COL[4003] = 1'b1;
assign COL[4004] = 1'b1;
assign COL[4005] = 1'b1;
assign COL[4006] = 1'b0;
assign COL[4007] = 1'b0;
assign COL[4008] = 1'b0;
assign COL[4009] = 1'b0;
assign COL[4010] = 1'b0;
assign COL[4011] = 1'b0;
assign COL[4012] = 1'b0;
assign COL[4013] = 1'b0;
assign COL[4014] = 1'b0;
assign COL[4015] = 1'b0;
assign COL[4016] = 1'b1;
assign COL[4017] = 1'b1;
assign COL[4018] = 1'b1;
assign COL[4019] = 1'b1;
assign COL[4020] = 1'b0;
assign COL[4021] = 1'b0;
assign COL[4022] = 1'b0;
assign COL[4023] = 1'b0;
assign COL[4024] = 1'b0;
assign COL[4025] = 1'b0;
assign COL[4026] = 1'b0;
assign COL[4027] = 1'b0;
assign COL[4028] = 1'b0;
assign COL[4029] = 1'b0;
assign COL[4030] = 1'b0;
assign COL[4031] = 1'b0;
assign COL[4032] = 1'b0;
assign COL[4033] = 1'b0;
assign COL[4034] = 1'b0;
assign COL[4035] = 1'b0;
assign COL[4036] = 1'b0;
assign COL[4037] = 1'b0;
assign COL[4038] = 1'b0;
assign COL[4039] = 1'b0;
assign COL[4040] = 1'b1;
assign COL[4041] = 1'b1;
assign COL[4042] = 1'b1;
assign COL[4043] = 1'b1;
assign COL[4044] = 1'b0;
assign COL[4045] = 1'b0;
assign COL[4046] = 1'b0;
assign COL[4047] = 1'b0;
assign COL[4048] = 1'b0;
assign COL[4049] = 1'b0;
assign COL[4050] = 1'b1;
assign COL[4051] = 1'b1;
assign COL[4052] = 1'b1;
assign COL[4053] = 1'b1;
assign COL[4054] = 1'b1;
assign COL[4055] = 1'b1;
assign COL[4056] = 1'b1;
assign COL[4057] = 1'b1;
assign COL[4058] = 1'b1;
assign COL[4059] = 1'b1;
assign COL[4060] = 1'b1;
assign COL[4061] = 1'b1;
assign COL[4062] = 1'b1;
assign COL[4063] = 1'b1;
assign COL[4064] = 1'b1;
assign COL[4065] = 1'b1;
assign COL[4066] = 1'b0;
assign COL[4067] = 1'b0;
assign COL[4068] = 1'b0;
assign COL[4069] = 1'b0;
assign COL[4070] = 1'b0;
assign COL[4071] = 1'b0;
assign COL[4072] = 1'b0;
assign COL[4073] = 1'b0;
assign COL[4074] = 1'b0;
assign COL[4075] = 1'b0;
assign COL[4076] = 1'b0;
assign COL[4077] = 1'b0;
assign COL[4078] = 1'b0;
assign COL[4079] = 1'b0;
assign COL[4080] = 1'b0;
assign COL[4081] = 1'b0;
assign COL[4082] = 1'b0;
assign COL[4083] = 1'b0;
assign COL[4084] = 1'b0;
assign COL[4085] = 1'b0;
assign COL[4086] = 1'b0;
assign COL[4087] = 1'b0;
assign COL[4088] = 1'b0;
assign COL[4089] = 1'b0;
assign COL[4090] = 1'b1;
assign COL[4091] = 1'b1;
assign COL[4092] = 1'b1;
assign COL[4093] = 1'b1;
assign COL[4094] = 1'b1;
assign COL[4095] = 1'b0;
assign COL[4096] = 1'b0;
assign COL[4097] = 1'b0;
assign COL[4098] = 1'b0;
assign COL[4099] = 1'b0;
assign COL[4100] = 1'b0;
assign COL[4101] = 1'b0;
assign COL[4102] = 1'b0;
assign COL[4103] = 1'b0;
assign COL[4104] = 1'b0;
assign COL[4105] = 1'b0;
assign COL[4106] = 1'b0;
assign COL[4107] = 1'b0;
assign COL[4108] = 1'b0;
assign COL[4109] = 1'b0;
assign COL[4110] = 1'b0;
assign COL[4111] = 1'b0;
assign COL[4112] = 1'b0;
assign COL[4113] = 1'b0;
assign COL[4114] = 1'b0;
assign COL[4115] = 1'b0;
assign COL[4116] = 1'b0;
assign COL[4117] = 1'b0;
assign COL[4118] = 1'b0;
assign COL[4119] = 1'b0;
assign COL[4120] = 1'b0;
assign COL[4121] = 1'b0;
assign COL[4122] = 1'b0;
assign COL[4123] = 1'b0;
assign COL[4124] = 1'b0;
assign COL[4125] = 1'b0;
assign COL[4126] = 1'b0;
assign COL[4127] = 1'b0;
assign COL[4128] = 1'b0;
assign COL[4129] = 1'b0;
assign COL[4130] = 1'b0;
assign COL[4131] = 1'b0;
assign COL[4132] = 1'b0;
assign COL[4133] = 1'b0;
assign COL[4134] = 1'b0;
assign COL[4135] = 1'b0;
assign COL[4136] = 1'b0;
assign COL[4137] = 1'b0;
assign COL[4138] = 1'b0;
assign COL[4139] = 1'b0;
assign COL[4140] = 1'b0;
assign COL[4141] = 1'b0;
assign COL[4142] = 1'b0;
assign COL[4143] = 1'b0;
assign COL[4144] = 1'b0;
assign COL[4145] = 1'b0;
assign COL[4146] = 1'b0;
assign COL[4147] = 1'b0;
assign COL[4148] = 1'b0;
assign COL[4149] = 1'b0;
assign COL[4150] = 1'b0;
assign COL[4151] = 1'b0;
assign COL[4152] = 1'b0;
assign COL[4153] = 1'b0;
assign COL[4154] = 1'b0;
assign COL[4155] = 1'b0;
assign COL[4156] = 1'b0;
assign COL[4157] = 1'b0;
assign COL[4158] = 1'b0;
assign COL[4159] = 1'b0;
assign COL[4160] = 1'b0;
assign COL[4161] = 1'b1;
assign COL[4162] = 1'b1;
assign COL[4163] = 1'b1;
assign COL[4164] = 1'b1;
assign COL[4165] = 1'b1;
assign COL[4166] = 1'b0;
assign COL[4167] = 1'b0;
assign COL[4168] = 1'b0;
assign COL[4169] = 1'b0;
assign COL[4170] = 1'b0;
assign COL[4171] = 1'b0;
assign COL[4172] = 1'b0;
assign COL[4173] = 1'b0;
assign COL[4174] = 1'b0;
assign COL[4175] = 1'b0;
assign COL[4176] = 1'b1;
assign COL[4177] = 1'b1;
assign COL[4178] = 1'b1;
assign COL[4179] = 1'b1;
assign COL[4180] = 1'b0;
assign COL[4181] = 1'b0;
assign COL[4182] = 1'b0;
assign COL[4183] = 1'b0;
assign COL[4184] = 1'b0;
assign COL[4185] = 1'b0;
assign COL[4186] = 1'b0;
assign COL[4187] = 1'b0;
assign COL[4188] = 1'b0;
assign COL[4189] = 1'b0;
assign COL[4190] = 1'b0;
assign COL[4191] = 1'b0;
assign COL[4192] = 1'b0;
assign COL[4193] = 1'b0;
assign COL[4194] = 1'b0;
assign COL[4195] = 1'b0;
assign COL[4196] = 1'b0;
assign COL[4197] = 1'b0;
assign COL[4198] = 1'b0;
assign COL[4199] = 1'b0;
assign COL[4200] = 1'b1;
assign COL[4201] = 1'b1;
assign COL[4202] = 1'b1;
assign COL[4203] = 1'b1;
assign COL[4204] = 1'b0;
assign COL[4205] = 1'b0;
assign COL[4206] = 1'b0;
assign COL[4207] = 1'b0;
assign COL[4208] = 1'b0;
assign COL[4209] = 1'b0;
assign COL[4210] = 1'b1;
assign COL[4211] = 1'b1;
assign COL[4212] = 1'b1;
assign COL[4213] = 1'b1;
assign COL[4214] = 1'b1;
assign COL[4215] = 1'b1;
assign COL[4216] = 1'b1;
assign COL[4217] = 1'b1;
assign COL[4218] = 1'b1;
assign COL[4219] = 1'b1;
assign COL[4220] = 1'b1;
assign COL[4221] = 1'b1;
assign COL[4222] = 1'b1;
assign COL[4223] = 1'b1;
assign COL[4224] = 1'b1;
assign COL[4225] = 1'b1;
assign COL[4226] = 1'b0;
assign COL[4227] = 1'b0;
assign COL[4228] = 1'b0;
assign COL[4229] = 1'b0;
assign COL[4230] = 1'b0;
assign COL[4231] = 1'b0;
assign COL[4232] = 1'b0;
assign COL[4233] = 1'b0;
assign COL[4234] = 1'b0;
assign COL[4235] = 1'b0;
assign COL[4236] = 1'b0;
assign COL[4237] = 1'b0;
assign COL[4238] = 1'b0;
assign COL[4239] = 1'b0;
assign COL[4240] = 1'b0;
assign COL[4241] = 1'b0;
assign COL[4242] = 1'b0;
assign COL[4243] = 1'b0;
assign COL[4244] = 1'b0;
assign COL[4245] = 1'b0;
assign COL[4246] = 1'b0;
assign COL[4247] = 1'b0;
assign COL[4248] = 1'b0;
assign COL[4249] = 1'b0;
assign COL[4250] = 1'b1;
assign COL[4251] = 1'b1;
assign COL[4252] = 1'b1;
assign COL[4253] = 1'b1;
assign COL[4254] = 1'b1;
assign COL[4255] = 1'b0;
assign COL[4256] = 1'b0;
assign COL[4257] = 1'b0;
assign COL[4258] = 1'b0;
assign COL[4259] = 1'b0;
assign COL[4260] = 1'b0;
assign COL[4261] = 1'b0;
assign COL[4262] = 1'b0;
assign COL[4263] = 1'b0;
assign COL[4264] = 1'b0;
assign COL[4265] = 1'b0;
assign COL[4266] = 1'b0;
assign COL[4267] = 1'b0;
assign COL[4268] = 1'b0;
assign COL[4269] = 1'b0;
assign COL[4270] = 1'b0;
assign COL[4271] = 1'b0;
assign COL[4272] = 1'b0;
assign COL[4273] = 1'b0;
assign COL[4274] = 1'b0;
assign COL[4275] = 1'b0;
assign COL[4276] = 1'b0;
assign COL[4277] = 1'b0;
assign COL[4278] = 1'b0;
assign COL[4279] = 1'b0;
assign COL[4280] = 1'b0;
assign COL[4281] = 1'b0;
assign COL[4282] = 1'b0;
assign COL[4283] = 1'b0;
assign COL[4284] = 1'b0;
assign COL[4285] = 1'b0;
assign COL[4286] = 1'b0;
assign COL[4287] = 1'b0;
assign COL[4288] = 1'b0;
assign COL[4289] = 1'b0;
assign COL[4290] = 1'b0;
assign COL[4291] = 1'b0;
assign COL[4292] = 1'b0;
assign COL[4293] = 1'b0;
assign COL[4294] = 1'b0;
assign COL[4295] = 1'b0;
assign COL[4296] = 1'b0;
assign COL[4297] = 1'b0;
assign COL[4298] = 1'b0;
assign COL[4299] = 1'b0;
assign COL[4300] = 1'b0;
assign COL[4301] = 1'b0;
assign COL[4302] = 1'b0;
assign COL[4303] = 1'b0;
assign COL[4304] = 1'b0;
assign COL[4305] = 1'b0;
assign COL[4306] = 1'b0;
assign COL[4307] = 1'b0;
assign COL[4308] = 1'b0;
assign COL[4309] = 1'b0;
assign COL[4310] = 1'b0;
assign COL[4311] = 1'b0;
assign COL[4312] = 1'b0;
assign COL[4313] = 1'b0;
assign COL[4314] = 1'b0;
assign COL[4315] = 1'b0;
assign COL[4316] = 1'b0;
assign COL[4317] = 1'b0;
assign COL[4318] = 1'b0;
assign COL[4319] = 1'b0;
assign COL[4320] = 1'b0;
assign COL[4321] = 1'b1;
assign COL[4322] = 1'b1;
assign COL[4323] = 1'b1;
assign COL[4324] = 1'b1;
assign COL[4325] = 1'b1;
assign COL[4326] = 1'b0;
assign COL[4327] = 1'b0;
assign COL[4328] = 1'b0;
assign COL[4329] = 1'b0;
assign COL[4330] = 1'b0;
assign COL[4331] = 1'b0;
assign COL[4332] = 1'b0;
assign COL[4333] = 1'b0;
assign COL[4334] = 1'b0;
assign COL[4335] = 1'b0;
assign COL[4336] = 1'b1;
assign COL[4337] = 1'b1;
assign COL[4338] = 1'b1;
assign COL[4339] = 1'b1;
assign COL[4340] = 1'b0;
assign COL[4341] = 1'b0;
assign COL[4342] = 1'b0;
assign COL[4343] = 1'b0;
assign COL[4344] = 1'b0;
assign COL[4345] = 1'b0;
assign COL[4346] = 1'b0;
assign COL[4347] = 1'b0;
assign COL[4348] = 1'b0;
assign COL[4349] = 1'b0;
assign COL[4350] = 1'b0;
assign COL[4351] = 1'b0;
assign COL[4352] = 1'b0;
assign COL[4353] = 1'b0;
assign COL[4354] = 1'b0;
assign COL[4355] = 1'b0;
assign COL[4356] = 1'b0;
assign COL[4357] = 1'b0;
assign COL[4358] = 1'b0;
assign COL[4359] = 1'b0;
assign COL[4360] = 1'b1;
assign COL[4361] = 1'b1;
assign COL[4362] = 1'b1;
assign COL[4363] = 1'b1;
assign COL[4364] = 1'b0;
assign COL[4365] = 1'b0;
assign COL[4366] = 1'b0;
assign COL[4367] = 1'b0;
assign COL[4368] = 1'b0;
assign COL[4369] = 1'b0;
assign COL[4370] = 1'b0;
assign COL[4371] = 1'b0;
assign COL[4372] = 1'b0;
assign COL[4373] = 1'b0;
assign COL[4374] = 1'b0;
assign COL[4375] = 1'b0;
assign COL[4376] = 1'b0;
assign COL[4377] = 1'b0;
assign COL[4378] = 1'b0;
assign COL[4379] = 1'b0;
assign COL[4380] = 1'b0;
assign COL[4381] = 1'b1;
assign COL[4382] = 1'b1;
assign COL[4383] = 1'b1;
assign COL[4384] = 1'b1;
assign COL[4385] = 1'b1;
assign COL[4386] = 1'b0;
assign COL[4387] = 1'b0;
assign COL[4388] = 1'b0;
assign COL[4389] = 1'b0;
assign COL[4390] = 1'b0;
assign COL[4391] = 1'b0;
assign COL[4392] = 1'b0;
assign COL[4393] = 1'b0;
assign COL[4394] = 1'b0;
assign COL[4395] = 1'b0;
assign COL[4396] = 1'b0;
assign COL[4397] = 1'b0;
assign COL[4398] = 1'b0;
assign COL[4399] = 1'b0;
assign COL[4400] = 1'b0;
assign COL[4401] = 1'b0;
assign COL[4402] = 1'b0;
assign COL[4403] = 1'b0;
assign COL[4404] = 1'b0;
assign COL[4405] = 1'b0;
assign COL[4406] = 1'b0;
assign COL[4407] = 1'b0;
assign COL[4408] = 1'b0;
assign COL[4409] = 1'b0;
assign COL[4410] = 1'b1;
assign COL[4411] = 1'b1;
assign COL[4412] = 1'b1;
assign COL[4413] = 1'b1;
assign COL[4414] = 1'b1;
assign COL[4415] = 1'b0;
assign COL[4416] = 1'b0;
assign COL[4417] = 1'b0;
assign COL[4418] = 1'b0;
assign COL[4419] = 1'b0;
assign COL[4420] = 1'b0;
assign COL[4421] = 1'b0;
assign COL[4422] = 1'b0;
assign COL[4423] = 1'b0;
assign COL[4424] = 1'b0;
assign COL[4425] = 1'b0;
assign COL[4426] = 1'b0;
assign COL[4427] = 1'b0;
assign COL[4428] = 1'b0;
assign COL[4429] = 1'b0;
assign COL[4430] = 1'b0;
assign COL[4431] = 1'b0;
assign COL[4432] = 1'b0;
assign COL[4433] = 1'b0;
assign COL[4434] = 1'b0;
assign COL[4435] = 1'b0;
assign COL[4436] = 1'b0;
assign COL[4437] = 1'b0;
assign COL[4438] = 1'b0;
assign COL[4439] = 1'b0;
assign COL[4440] = 1'b0;
assign COL[4441] = 1'b0;
assign COL[4442] = 1'b0;
assign COL[4443] = 1'b0;
assign COL[4444] = 1'b0;
assign COL[4445] = 1'b0;
assign COL[4446] = 1'b0;
assign COL[4447] = 1'b0;
assign COL[4448] = 1'b0;
assign COL[4449] = 1'b0;
assign COL[4450] = 1'b0;
assign COL[4451] = 1'b0;
assign COL[4452] = 1'b0;
assign COL[4453] = 1'b0;
assign COL[4454] = 1'b0;
assign COL[4455] = 1'b0;
assign COL[4456] = 1'b0;
assign COL[4457] = 1'b0;
assign COL[4458] = 1'b0;
assign COL[4459] = 1'b0;
assign COL[4460] = 1'b0;
assign COL[4461] = 1'b0;
assign COL[4462] = 1'b0;
assign COL[4463] = 1'b0;
assign COL[4464] = 1'b0;
assign COL[4465] = 1'b0;
assign COL[4466] = 1'b0;
assign COL[4467] = 1'b0;
assign COL[4468] = 1'b0;
assign COL[4469] = 1'b0;
assign COL[4470] = 1'b0;
assign COL[4471] = 1'b0;
assign COL[4472] = 1'b0;
assign COL[4473] = 1'b0;
assign COL[4474] = 1'b0;
assign COL[4475] = 1'b0;
assign COL[4476] = 1'b0;
assign COL[4477] = 1'b0;
assign COL[4478] = 1'b0;
assign COL[4479] = 1'b0;
assign COL[4480] = 1'b0;
assign COL[4481] = 1'b1;
assign COL[4482] = 1'b1;
assign COL[4483] = 1'b1;
assign COL[4484] = 1'b1;
assign COL[4485] = 1'b1;
assign COL[4486] = 1'b0;
assign COL[4487] = 1'b0;
assign COL[4488] = 1'b0;
assign COL[4489] = 1'b0;
assign COL[4490] = 1'b0;
assign COL[4491] = 1'b0;
assign COL[4492] = 1'b0;
assign COL[4493] = 1'b0;
assign COL[4494] = 1'b0;
assign COL[4495] = 1'b0;
assign COL[4496] = 1'b1;
assign COL[4497] = 1'b1;
assign COL[4498] = 1'b1;
assign COL[4499] = 1'b1;
assign COL[4500] = 1'b0;
assign COL[4501] = 1'b0;
assign COL[4502] = 1'b0;
assign COL[4503] = 1'b0;
assign COL[4504] = 1'b0;
assign COL[4505] = 1'b0;
assign COL[4506] = 1'b0;
assign COL[4507] = 1'b0;
assign COL[4508] = 1'b0;
assign COL[4509] = 1'b0;
assign COL[4510] = 1'b0;
assign COL[4511] = 1'b0;
assign COL[4512] = 1'b0;
assign COL[4513] = 1'b0;
assign COL[4514] = 1'b0;
assign COL[4515] = 1'b0;
assign COL[4516] = 1'b0;
assign COL[4517] = 1'b0;
assign COL[4518] = 1'b0;
assign COL[4519] = 1'b0;
assign COL[4520] = 1'b1;
assign COL[4521] = 1'b1;
assign COL[4522] = 1'b1;
assign COL[4523] = 1'b1;
assign COL[4524] = 1'b0;
assign COL[4525] = 1'b0;
assign COL[4526] = 1'b0;
assign COL[4527] = 1'b0;
assign COL[4528] = 1'b0;
assign COL[4529] = 1'b0;
assign COL[4530] = 1'b0;
assign COL[4531] = 1'b0;
assign COL[4532] = 1'b0;
assign COL[4533] = 1'b0;
assign COL[4534] = 1'b0;
assign COL[4535] = 1'b0;
assign COL[4536] = 1'b0;
assign COL[4537] = 1'b0;
assign COL[4538] = 1'b0;
assign COL[4539] = 1'b0;
assign COL[4540] = 1'b0;
assign COL[4541] = 1'b1;
assign COL[4542] = 1'b1;
assign COL[4543] = 1'b1;
assign COL[4544] = 1'b1;
assign COL[4545] = 1'b1;
assign COL[4546] = 1'b0;
assign COL[4547] = 1'b0;
assign COL[4548] = 1'b0;
assign COL[4549] = 1'b0;
assign COL[4550] = 1'b0;
assign COL[4551] = 1'b0;
assign COL[4552] = 1'b0;
assign COL[4553] = 1'b0;
assign COL[4554] = 1'b0;
assign COL[4555] = 1'b0;
assign COL[4556] = 1'b0;
assign COL[4557] = 1'b0;
assign COL[4558] = 1'b0;
assign COL[4559] = 1'b0;
assign COL[4560] = 1'b0;
assign COL[4561] = 1'b0;
assign COL[4562] = 1'b0;
assign COL[4563] = 1'b0;
assign COL[4564] = 1'b0;
assign COL[4565] = 1'b0;
assign COL[4566] = 1'b0;
assign COL[4567] = 1'b0;
assign COL[4568] = 1'b0;
assign COL[4569] = 1'b0;
assign COL[4570] = 1'b1;
assign COL[4571] = 1'b1;
assign COL[4572] = 1'b1;
assign COL[4573] = 1'b1;
assign COL[4574] = 1'b1;
assign COL[4575] = 1'b0;
assign COL[4576] = 1'b0;
assign COL[4577] = 1'b0;
assign COL[4578] = 1'b0;
assign COL[4579] = 1'b0;
assign COL[4580] = 1'b0;
assign COL[4581] = 1'b0;
assign COL[4582] = 1'b0;
assign COL[4583] = 1'b0;
assign COL[4584] = 1'b0;
assign COL[4585] = 1'b0;
assign COL[4586] = 1'b0;
assign COL[4587] = 1'b0;
assign COL[4588] = 1'b0;
assign COL[4589] = 1'b0;
assign COL[4590] = 1'b0;
assign COL[4591] = 1'b0;
assign COL[4592] = 1'b0;
assign COL[4593] = 1'b0;
assign COL[4594] = 1'b0;
assign COL[4595] = 1'b0;
assign COL[4596] = 1'b0;
assign COL[4597] = 1'b0;
assign COL[4598] = 1'b0;
assign COL[4599] = 1'b0;
assign COL[4600] = 1'b0;
assign COL[4601] = 1'b0;
assign COL[4602] = 1'b0;
assign COL[4603] = 1'b0;
assign COL[4604] = 1'b0;
assign COL[4605] = 1'b0;
assign COL[4606] = 1'b0;
assign COL[4607] = 1'b0;
assign COL[4608] = 1'b0;
assign COL[4609] = 1'b0;
assign COL[4610] = 1'b0;
assign COL[4611] = 1'b0;
assign COL[4612] = 1'b0;
assign COL[4613] = 1'b0;
assign COL[4614] = 1'b0;
assign COL[4615] = 1'b0;
assign COL[4616] = 1'b0;
assign COL[4617] = 1'b0;
assign COL[4618] = 1'b0;
assign COL[4619] = 1'b0;
assign COL[4620] = 1'b0;
assign COL[4621] = 1'b0;
assign COL[4622] = 1'b0;
assign COL[4623] = 1'b0;
assign COL[4624] = 1'b0;
assign COL[4625] = 1'b0;
assign COL[4626] = 1'b0;
assign COL[4627] = 1'b0;
assign COL[4628] = 1'b0;
assign COL[4629] = 1'b0;
assign COL[4630] = 1'b0;
assign COL[4631] = 1'b0;
assign COL[4632] = 1'b0;
assign COL[4633] = 1'b0;
assign COL[4634] = 1'b0;
assign COL[4635] = 1'b0;
assign COL[4636] = 1'b0;
assign COL[4637] = 1'b0;
assign COL[4638] = 1'b0;
assign COL[4639] = 1'b0;
assign COL[4640] = 1'b0;
assign COL[4641] = 1'b1;
assign COL[4642] = 1'b1;
assign COL[4643] = 1'b1;
assign COL[4644] = 1'b1;
assign COL[4645] = 1'b1;
assign COL[4646] = 1'b0;
assign COL[4647] = 1'b0;
assign COL[4648] = 1'b0;
assign COL[4649] = 1'b0;
assign COL[4650] = 1'b0;
assign COL[4651] = 1'b0;
assign COL[4652] = 1'b0;
assign COL[4653] = 1'b0;
assign COL[4654] = 1'b0;
assign COL[4655] = 1'b0;
assign COL[4656] = 1'b1;
assign COL[4657] = 1'b1;
assign COL[4658] = 1'b1;
assign COL[4659] = 1'b1;
assign COL[4660] = 1'b0;
assign COL[4661] = 1'b0;
assign COL[4662] = 1'b0;
assign COL[4663] = 1'b0;
assign COL[4664] = 1'b0;
assign COL[4665] = 1'b0;
assign COL[4666] = 1'b0;
assign COL[4667] = 1'b0;
assign COL[4668] = 1'b0;
assign COL[4669] = 1'b0;
assign COL[4670] = 1'b0;
assign COL[4671] = 1'b0;
assign COL[4672] = 1'b0;
assign COL[4673] = 1'b0;
assign COL[4674] = 1'b0;
assign COL[4675] = 1'b0;
assign COL[4676] = 1'b0;
assign COL[4677] = 1'b0;
assign COL[4678] = 1'b0;
assign COL[4679] = 1'b0;
assign COL[4680] = 1'b1;
assign COL[4681] = 1'b1;
assign COL[4682] = 1'b1;
assign COL[4683] = 1'b1;
assign COL[4684] = 1'b0;
assign COL[4685] = 1'b0;
assign COL[4686] = 1'b0;
assign COL[4687] = 1'b0;
assign COL[4688] = 1'b0;
assign COL[4689] = 1'b0;
assign COL[4690] = 1'b0;
assign COL[4691] = 1'b0;
assign COL[4692] = 1'b0;
assign COL[4693] = 1'b0;
assign COL[4694] = 1'b0;
assign COL[4695] = 1'b0;
assign COL[4696] = 1'b0;
assign COL[4697] = 1'b0;
assign COL[4698] = 1'b0;
assign COL[4699] = 1'b0;
assign COL[4700] = 1'b0;
assign COL[4701] = 1'b1;
assign COL[4702] = 1'b1;
assign COL[4703] = 1'b1;
assign COL[4704] = 1'b1;
assign COL[4705] = 1'b1;
assign COL[4706] = 1'b0;
assign COL[4707] = 1'b0;
assign COL[4708] = 1'b0;
assign COL[4709] = 1'b0;
assign COL[4710] = 1'b0;
assign COL[4711] = 1'b0;
assign COL[4712] = 1'b0;
assign COL[4713] = 1'b0;
assign COL[4714] = 1'b0;
assign COL[4715] = 1'b0;
assign COL[4716] = 1'b0;
assign COL[4717] = 1'b0;
assign COL[4718] = 1'b0;
assign COL[4719] = 1'b0;
assign COL[4720] = 1'b0;
assign COL[4721] = 1'b0;
assign COL[4722] = 1'b0;
assign COL[4723] = 1'b0;
assign COL[4724] = 1'b0;
assign COL[4725] = 1'b0;
assign COL[4726] = 1'b0;
assign COL[4727] = 1'b0;
assign COL[4728] = 1'b0;
assign COL[4729] = 1'b0;
assign COL[4730] = 1'b1;
assign COL[4731] = 1'b1;
assign COL[4732] = 1'b1;
assign COL[4733] = 1'b1;
assign COL[4734] = 1'b1;
assign COL[4735] = 1'b0;
assign COL[4736] = 1'b0;
assign COL[4737] = 1'b0;
assign COL[4738] = 1'b0;
assign COL[4739] = 1'b0;
assign COL[4740] = 1'b0;
assign COL[4741] = 1'b0;
assign COL[4742] = 1'b0;
assign COL[4743] = 1'b0;
assign COL[4744] = 1'b0;
assign COL[4745] = 1'b0;
assign COL[4746] = 1'b0;
assign COL[4747] = 1'b0;
assign COL[4748] = 1'b0;
assign COL[4749] = 1'b0;
assign COL[4750] = 1'b0;
assign COL[4751] = 1'b0;
assign COL[4752] = 1'b0;
assign COL[4753] = 1'b0;
assign COL[4754] = 1'b0;
assign COL[4755] = 1'b0;
assign COL[4756] = 1'b0;
assign COL[4757] = 1'b0;
assign COL[4758] = 1'b0;
assign COL[4759] = 1'b0;
assign COL[4760] = 1'b0;
assign COL[4761] = 1'b0;
assign COL[4762] = 1'b0;
assign COL[4763] = 1'b0;
assign COL[4764] = 1'b0;
assign COL[4765] = 1'b0;
assign COL[4766] = 1'b0;
assign COL[4767] = 1'b0;
assign COL[4768] = 1'b0;
assign COL[4769] = 1'b0;
assign COL[4770] = 1'b0;
assign COL[4771] = 1'b0;
assign COL[4772] = 1'b0;
assign COL[4773] = 1'b0;
assign COL[4774] = 1'b0;
assign COL[4775] = 1'b0;
assign COL[4776] = 1'b0;
assign COL[4777] = 1'b0;
assign COL[4778] = 1'b0;
assign COL[4779] = 1'b0;
assign COL[4780] = 1'b0;
assign COL[4781] = 1'b0;
assign COL[4782] = 1'b0;
assign COL[4783] = 1'b0;
assign COL[4784] = 1'b0;
assign COL[4785] = 1'b0;
assign COL[4786] = 1'b0;
assign COL[4787] = 1'b0;
assign COL[4788] = 1'b0;
assign COL[4789] = 1'b0;
assign COL[4790] = 1'b0;
assign COL[4791] = 1'b0;
assign COL[4792] = 1'b0;
assign COL[4793] = 1'b0;
assign COL[4794] = 1'b0;
assign COL[4795] = 1'b0;
assign COL[4796] = 1'b0;
assign COL[4797] = 1'b0;
assign COL[4798] = 1'b0;
assign COL[4799] = 1'b0;
assign COL[4800] = 1'b0;
assign COL[4801] = 1'b1;
assign COL[4802] = 1'b1;
assign COL[4803] = 1'b1;
assign COL[4804] = 1'b1;
assign COL[4805] = 1'b1;
assign COL[4806] = 1'b0;
assign COL[4807] = 1'b0;
assign COL[4808] = 1'b0;
assign COL[4809] = 1'b0;
assign COL[4810] = 1'b0;
assign COL[4811] = 1'b0;
assign COL[4812] = 1'b0;
assign COL[4813] = 1'b0;
assign COL[4814] = 1'b0;
assign COL[4815] = 1'b0;
assign COL[4816] = 1'b1;
assign COL[4817] = 1'b1;
assign COL[4818] = 1'b1;
assign COL[4819] = 1'b1;
assign COL[4820] = 1'b0;
assign COL[4821] = 1'b0;
assign COL[4822] = 1'b0;
assign COL[4823] = 1'b0;
assign COL[4824] = 1'b0;
assign COL[4825] = 1'b0;
assign COL[4826] = 1'b0;
assign COL[4827] = 1'b0;
assign COL[4828] = 1'b0;
assign COL[4829] = 1'b0;
assign COL[4830] = 1'b0;
assign COL[4831] = 1'b0;
assign COL[4832] = 1'b0;
assign COL[4833] = 1'b0;
assign COL[4834] = 1'b0;
assign COL[4835] = 1'b0;
assign COL[4836] = 1'b0;
assign COL[4837] = 1'b0;
assign COL[4838] = 1'b0;
assign COL[4839] = 1'b0;
assign COL[4840] = 1'b1;
assign COL[4841] = 1'b1;
assign COL[4842] = 1'b1;
assign COL[4843] = 1'b1;
assign COL[4844] = 1'b0;
assign COL[4845] = 1'b0;
assign COL[4846] = 1'b0;
assign COL[4847] = 1'b0;
assign COL[4848] = 1'b0;
assign COL[4849] = 1'b0;
assign COL[4850] = 1'b0;
assign COL[4851] = 1'b0;
assign COL[4852] = 1'b0;
assign COL[4853] = 1'b0;
assign COL[4854] = 1'b0;
assign COL[4855] = 1'b0;
assign COL[4856] = 1'b0;
assign COL[4857] = 1'b0;
assign COL[4858] = 1'b0;
assign COL[4859] = 1'b0;
assign COL[4860] = 1'b0;
assign COL[4861] = 1'b1;
assign COL[4862] = 1'b1;
assign COL[4863] = 1'b1;
assign COL[4864] = 1'b1;
assign COL[4865] = 1'b1;
assign COL[4866] = 1'b0;
assign COL[4867] = 1'b0;
assign COL[4868] = 1'b0;
assign COL[4869] = 1'b0;
assign COL[4870] = 1'b0;
assign COL[4871] = 1'b0;
assign COL[4872] = 1'b0;
assign COL[4873] = 1'b0;
assign COL[4874] = 1'b0;
assign COL[4875] = 1'b0;
assign COL[4876] = 1'b0;
assign COL[4877] = 1'b0;
assign COL[4878] = 1'b0;
assign COL[4879] = 1'b0;
assign COL[4880] = 1'b0;
assign COL[4881] = 1'b0;
assign COL[4882] = 1'b0;
assign COL[4883] = 1'b0;
assign COL[4884] = 1'b0;
assign COL[4885] = 1'b0;
assign COL[4886] = 1'b0;
assign COL[4887] = 1'b0;
assign COL[4888] = 1'b0;
assign COL[4889] = 1'b0;
assign COL[4890] = 1'b1;
assign COL[4891] = 1'b1;
assign COL[4892] = 1'b1;
assign COL[4893] = 1'b1;
assign COL[4894] = 1'b1;
assign COL[4895] = 1'b0;
assign COL[4896] = 1'b0;
assign COL[4897] = 1'b0;
assign COL[4898] = 1'b0;
assign COL[4899] = 1'b0;
assign COL[4900] = 1'b0;
assign COL[4901] = 1'b0;
assign COL[4902] = 1'b0;
assign COL[4903] = 1'b0;
assign COL[4904] = 1'b0;
assign COL[4905] = 1'b0;
assign COL[4906] = 1'b0;
assign COL[4907] = 1'b0;
assign COL[4908] = 1'b0;
assign COL[4909] = 1'b0;
assign COL[4910] = 1'b0;
assign COL[4911] = 1'b0;
assign COL[4912] = 1'b0;
assign COL[4913] = 1'b0;
assign COL[4914] = 1'b0;
assign COL[4915] = 1'b0;
assign COL[4916] = 1'b0;
assign COL[4917] = 1'b0;
assign COL[4918] = 1'b0;
assign COL[4919] = 1'b0;
assign COL[4920] = 1'b0;
assign COL[4921] = 1'b0;
assign COL[4922] = 1'b0;
assign COL[4923] = 1'b0;
assign COL[4924] = 1'b0;
assign COL[4925] = 1'b0;
assign COL[4926] = 1'b0;
assign COL[4927] = 1'b0;
assign COL[4928] = 1'b0;
assign COL[4929] = 1'b0;
assign COL[4930] = 1'b0;
assign COL[4931] = 1'b0;
assign COL[4932] = 1'b0;
assign COL[4933] = 1'b0;
assign COL[4934] = 1'b0;
assign COL[4935] = 1'b0;
assign COL[4936] = 1'b0;
assign COL[4937] = 1'b0;
assign COL[4938] = 1'b0;
assign COL[4939] = 1'b0;
assign COL[4940] = 1'b0;
assign COL[4941] = 1'b0;
assign COL[4942] = 1'b0;
assign COL[4943] = 1'b0;
assign COL[4944] = 1'b0;
assign COL[4945] = 1'b0;
assign COL[4946] = 1'b0;
assign COL[4947] = 1'b0;
assign COL[4948] = 1'b0;
assign COL[4949] = 1'b0;
assign COL[4950] = 1'b0;
assign COL[4951] = 1'b0;
assign COL[4952] = 1'b0;
assign COL[4953] = 1'b0;
assign COL[4954] = 1'b0;
assign COL[4955] = 1'b0;
assign COL[4956] = 1'b0;
assign COL[4957] = 1'b0;
assign COL[4958] = 1'b0;
assign COL[4959] = 1'b0;
assign COL[4960] = 1'b0;
assign COL[4961] = 1'b1;
assign COL[4962] = 1'b1;
assign COL[4963] = 1'b1;
assign COL[4964] = 1'b1;
assign COL[4965] = 1'b1;
assign COL[4966] = 1'b0;
assign COL[4967] = 1'b0;
assign COL[4968] = 1'b0;
assign COL[4969] = 1'b0;
assign COL[4970] = 1'b0;
assign COL[4971] = 1'b0;
assign COL[4972] = 1'b0;
assign COL[4973] = 1'b0;
assign COL[4974] = 1'b0;
assign COL[4975] = 1'b0;
assign COL[4976] = 1'b1;
assign COL[4977] = 1'b1;
assign COL[4978] = 1'b1;
assign COL[4979] = 1'b1;
assign COL[4980] = 1'b0;
assign COL[4981] = 1'b0;
assign COL[4982] = 1'b0;
assign COL[4983] = 1'b0;
assign COL[4984] = 1'b0;
assign COL[4985] = 1'b0;
assign COL[4986] = 1'b0;
assign COL[4987] = 1'b0;
assign COL[4988] = 1'b0;
assign COL[4989] = 1'b0;
assign COL[4990] = 1'b0;
assign COL[4991] = 1'b0;
assign COL[4992] = 1'b0;
assign COL[4993] = 1'b0;
assign COL[4994] = 1'b0;
assign COL[4995] = 1'b0;
assign COL[4996] = 1'b0;
assign COL[4997] = 1'b0;
assign COL[4998] = 1'b0;
assign COL[4999] = 1'b0;
assign COL[5000] = 1'b1;
assign COL[5001] = 1'b1;
assign COL[5002] = 1'b1;
assign COL[5003] = 1'b1;
assign COL[5004] = 1'b0;
assign COL[5005] = 1'b0;
assign COL[5006] = 1'b0;
assign COL[5007] = 1'b0;
assign COL[5008] = 1'b0;
assign COL[5009] = 1'b0;
assign COL[5010] = 1'b0;
assign COL[5011] = 1'b0;
assign COL[5012] = 1'b0;
assign COL[5013] = 1'b0;
assign COL[5014] = 1'b0;
assign COL[5015] = 1'b0;
assign COL[5016] = 1'b0;
assign COL[5017] = 1'b0;
assign COL[5018] = 1'b0;
assign COL[5019] = 1'b0;
assign COL[5020] = 1'b0;
assign COL[5021] = 1'b1;
assign COL[5022] = 1'b1;
assign COL[5023] = 1'b1;
assign COL[5024] = 1'b1;
assign COL[5025] = 1'b1;
assign COL[5026] = 1'b0;
assign COL[5027] = 1'b0;
assign COL[5028] = 1'b0;
assign COL[5029] = 1'b0;
assign COL[5030] = 1'b0;
assign COL[5031] = 1'b0;
assign COL[5032] = 1'b0;
assign COL[5033] = 1'b0;
assign COL[5034] = 1'b0;
assign COL[5035] = 1'b0;
assign COL[5036] = 1'b0;
assign COL[5037] = 1'b0;
assign COL[5038] = 1'b0;
assign COL[5039] = 1'b0;
assign COL[5040] = 1'b0;
assign COL[5041] = 1'b0;
assign COL[5042] = 1'b0;
assign COL[5043] = 1'b0;
assign COL[5044] = 1'b0;
assign COL[5045] = 1'b0;
assign COL[5046] = 1'b0;
assign COL[5047] = 1'b0;
assign COL[5048] = 1'b0;
assign COL[5049] = 1'b0;
assign COL[5050] = 1'b1;
assign COL[5051] = 1'b1;
assign COL[5052] = 1'b1;
assign COL[5053] = 1'b1;
assign COL[5054] = 1'b1;
assign COL[5055] = 1'b0;
assign COL[5056] = 1'b0;
assign COL[5057] = 1'b0;
assign COL[5058] = 1'b0;
assign COL[5059] = 1'b0;
assign COL[5060] = 1'b0;
assign COL[5061] = 1'b0;
assign COL[5062] = 1'b0;
assign COL[5063] = 1'b0;
assign COL[5064] = 1'b0;
assign COL[5065] = 1'b0;
assign COL[5066] = 1'b0;
assign COL[5067] = 1'b0;
assign COL[5068] = 1'b0;
assign COL[5069] = 1'b0;
assign COL[5070] = 1'b0;
assign COL[5071] = 1'b0;
assign COL[5072] = 1'b0;
assign COL[5073] = 1'b0;
assign COL[5074] = 1'b0;
assign COL[5075] = 1'b0;
assign COL[5076] = 1'b0;
assign COL[5077] = 1'b0;
assign COL[5078] = 1'b0;
assign COL[5079] = 1'b0;
assign COL[5080] = 1'b0;
assign COL[5081] = 1'b0;
assign COL[5082] = 1'b0;
assign COL[5083] = 1'b0;
assign COL[5084] = 1'b0;
assign COL[5085] = 1'b0;
assign COL[5086] = 1'b0;
assign COL[5087] = 1'b0;
assign COL[5088] = 1'b0;
assign COL[5089] = 1'b0;
assign COL[5090] = 1'b0;
assign COL[5091] = 1'b0;
assign COL[5092] = 1'b0;
assign COL[5093] = 1'b0;
assign COL[5094] = 1'b0;
assign COL[5095] = 1'b0;
assign COL[5096] = 1'b0;
assign COL[5097] = 1'b0;
assign COL[5098] = 1'b0;
assign COL[5099] = 1'b0;
assign COL[5100] = 1'b0;
assign COL[5101] = 1'b0;
assign COL[5102] = 1'b0;
assign COL[5103] = 1'b0;
assign COL[5104] = 1'b0;
assign COL[5105] = 1'b0;
assign COL[5106] = 1'b0;
assign COL[5107] = 1'b0;
assign COL[5108] = 1'b0;
assign COL[5109] = 1'b0;
assign COL[5110] = 1'b0;
assign COL[5111] = 1'b0;
assign COL[5112] = 1'b0;
assign COL[5113] = 1'b0;
assign COL[5114] = 1'b0;
assign COL[5115] = 1'b0;
assign COL[5116] = 1'b0;
assign COL[5117] = 1'b0;
assign COL[5118] = 1'b0;
assign COL[5119] = 1'b0;
assign COL[5120] = 1'b0;
assign COL[5121] = 1'b1;
assign COL[5122] = 1'b1;
assign COL[5123] = 1'b1;
assign COL[5124] = 1'b1;
assign COL[5125] = 1'b1;
assign COL[5126] = 1'b0;
assign COL[5127] = 1'b0;
assign COL[5128] = 1'b0;
assign COL[5129] = 1'b0;
assign COL[5130] = 1'b0;
assign COL[5131] = 1'b0;
assign COL[5132] = 1'b0;
assign COL[5133] = 1'b0;
assign COL[5134] = 1'b0;
assign COL[5135] = 1'b0;
assign COL[5136] = 1'b1;
assign COL[5137] = 1'b1;
assign COL[5138] = 1'b1;
assign COL[5139] = 1'b1;
assign COL[5140] = 1'b0;
assign COL[5141] = 1'b0;
assign COL[5142] = 1'b0;
assign COL[5143] = 1'b0;
assign COL[5144] = 1'b0;
assign COL[5145] = 1'b0;
assign COL[5146] = 1'b0;
assign COL[5147] = 1'b0;
assign COL[5148] = 1'b0;
assign COL[5149] = 1'b0;
assign COL[5150] = 1'b0;
assign COL[5151] = 1'b0;
assign COL[5152] = 1'b0;
assign COL[5153] = 1'b0;
assign COL[5154] = 1'b0;
assign COL[5155] = 1'b0;
assign COL[5156] = 1'b0;
assign COL[5157] = 1'b0;
assign COL[5158] = 1'b0;
assign COL[5159] = 1'b0;
assign COL[5160] = 1'b1;
assign COL[5161] = 1'b1;
assign COL[5162] = 1'b1;
assign COL[5163] = 1'b1;
assign COL[5164] = 1'b0;
assign COL[5165] = 1'b0;
assign COL[5166] = 1'b0;
assign COL[5167] = 1'b0;
assign COL[5168] = 1'b0;
assign COL[5169] = 1'b0;
assign COL[5170] = 1'b0;
assign COL[5171] = 1'b0;
assign COL[5172] = 1'b0;
assign COL[5173] = 1'b0;
assign COL[5174] = 1'b0;
assign COL[5175] = 1'b0;
assign COL[5176] = 1'b0;
assign COL[5177] = 1'b0;
assign COL[5178] = 1'b0;
assign COL[5179] = 1'b0;
assign COL[5180] = 1'b0;
assign COL[5181] = 1'b1;
assign COL[5182] = 1'b1;
assign COL[5183] = 1'b1;
assign COL[5184] = 1'b1;
assign COL[5185] = 1'b1;
assign COL[5186] = 1'b1;
assign COL[5187] = 1'b1;
assign COL[5188] = 1'b1;
assign COL[5189] = 1'b1;
assign COL[5190] = 1'b1;
assign COL[5191] = 1'b1;
assign COL[5192] = 1'b1;
assign COL[5193] = 1'b1;
assign COL[5194] = 1'b1;
assign COL[5195] = 1'b1;
assign COL[5196] = 1'b1;
assign COL[5197] = 1'b1;
assign COL[5198] = 1'b1;
assign COL[5199] = 1'b1;
assign COL[5200] = 1'b1;
assign COL[5201] = 1'b1;
assign COL[5202] = 1'b1;
assign COL[5203] = 1'b1;
assign COL[5204] = 1'b1;
assign COL[5205] = 1'b1;
assign COL[5206] = 1'b1;
assign COL[5207] = 1'b1;
assign COL[5208] = 1'b1;
assign COL[5209] = 1'b1;
assign COL[5210] = 1'b1;
assign COL[5211] = 1'b1;
assign COL[5212] = 1'b1;
assign COL[5213] = 1'b1;
assign COL[5214] = 1'b1;
assign COL[5215] = 1'b0;
assign COL[5216] = 1'b0;
assign COL[5217] = 1'b0;
assign COL[5218] = 1'b0;
assign COL[5219] = 1'b0;
assign COL[5220] = 1'b0;
assign COL[5221] = 1'b0;
assign COL[5222] = 1'b0;
assign COL[5223] = 1'b0;
assign COL[5224] = 1'b0;
assign COL[5225] = 1'b0;
assign COL[5226] = 1'b0;
assign COL[5227] = 1'b0;
assign COL[5228] = 1'b0;
assign COL[5229] = 1'b0;
assign COL[5230] = 1'b0;
assign COL[5231] = 1'b0;
assign COL[5232] = 1'b0;
assign COL[5233] = 1'b0;
assign COL[5234] = 1'b0;
assign COL[5235] = 1'b0;
assign COL[5236] = 1'b0;
assign COL[5237] = 1'b0;
assign COL[5238] = 1'b0;
assign COL[5239] = 1'b0;
assign COL[5240] = 1'b0;
assign COL[5241] = 1'b0;
assign COL[5242] = 1'b0;
assign COL[5243] = 1'b0;
assign COL[5244] = 1'b0;
assign COL[5245] = 1'b0;
assign COL[5246] = 1'b0;
assign COL[5247] = 1'b1;
assign COL[5248] = 1'b0;
assign COL[5249] = 1'b0;
assign COL[5250] = 1'b0;
assign COL[5251] = 1'b0;
assign COL[5252] = 1'b0;
assign COL[5253] = 1'b0;
assign COL[5254] = 1'b0;
assign COL[5255] = 1'b0;
assign COL[5256] = 1'b0;
assign COL[5257] = 1'b0;
assign COL[5258] = 1'b0;
assign COL[5259] = 1'b0;
assign COL[5260] = 1'b0;
assign COL[5261] = 1'b0;
assign COL[5262] = 1'b0;
assign COL[5263] = 1'b0;
assign COL[5264] = 1'b0;
assign COL[5265] = 1'b0;
assign COL[5266] = 1'b0;
assign COL[5267] = 1'b0;
assign COL[5268] = 1'b0;
assign COL[5269] = 1'b0;
assign COL[5270] = 1'b0;
assign COL[5271] = 1'b0;
assign COL[5272] = 1'b0;
assign COL[5273] = 1'b0;
assign COL[5274] = 1'b0;
assign COL[5275] = 1'b0;
assign COL[5276] = 1'b0;
assign COL[5277] = 1'b0;
assign COL[5278] = 1'b0;
assign COL[5279] = 1'b0;
assign COL[5280] = 1'b0;
assign COL[5281] = 1'b1;
assign COL[5282] = 1'b1;
assign COL[5283] = 1'b1;
assign COL[5284] = 1'b1;
assign COL[5285] = 1'b1;
assign COL[5286] = 1'b0;
assign COL[5287] = 1'b0;
assign COL[5288] = 1'b0;
assign COL[5289] = 1'b0;
assign COL[5290] = 1'b0;
assign COL[5291] = 1'b0;
assign COL[5292] = 1'b0;
assign COL[5293] = 1'b0;
assign COL[5294] = 1'b0;
assign COL[5295] = 1'b0;
assign COL[5296] = 1'b1;
assign COL[5297] = 1'b1;
assign COL[5298] = 1'b1;
assign COL[5299] = 1'b1;
assign COL[5300] = 1'b0;
assign COL[5301] = 1'b0;
assign COL[5302] = 1'b0;
assign COL[5303] = 1'b0;
assign COL[5304] = 1'b0;
assign COL[5305] = 1'b0;
assign COL[5306] = 1'b0;
assign COL[5307] = 1'b0;
assign COL[5308] = 1'b0;
assign COL[5309] = 1'b0;
assign COL[5310] = 1'b0;
assign COL[5311] = 1'b0;
assign COL[5312] = 1'b0;
assign COL[5313] = 1'b0;
assign COL[5314] = 1'b0;
assign COL[5315] = 1'b0;
assign COL[5316] = 1'b0;
assign COL[5317] = 1'b0;
assign COL[5318] = 1'b0;
assign COL[5319] = 1'b0;
assign COL[5320] = 1'b1;
assign COL[5321] = 1'b1;
assign COL[5322] = 1'b1;
assign COL[5323] = 1'b1;
assign COL[5324] = 1'b0;
assign COL[5325] = 1'b0;
assign COL[5326] = 1'b0;
assign COL[5327] = 1'b0;
assign COL[5328] = 1'b0;
assign COL[5329] = 1'b0;
assign COL[5330] = 1'b0;
assign COL[5331] = 1'b0;
assign COL[5332] = 1'b0;
assign COL[5333] = 1'b0;
assign COL[5334] = 1'b0;
assign COL[5335] = 1'b0;
assign COL[5336] = 1'b0;
assign COL[5337] = 1'b0;
assign COL[5338] = 1'b0;
assign COL[5339] = 1'b0;
assign COL[5340] = 1'b0;
assign COL[5341] = 1'b1;
assign COL[5342] = 1'b1;
assign COL[5343] = 1'b1;
assign COL[5344] = 1'b1;
assign COL[5345] = 1'b1;
assign COL[5346] = 1'b1;
assign COL[5347] = 1'b1;
assign COL[5348] = 1'b1;
assign COL[5349] = 1'b1;
assign COL[5350] = 1'b1;
assign COL[5351] = 1'b1;
assign COL[5352] = 1'b1;
assign COL[5353] = 1'b1;
assign COL[5354] = 1'b1;
assign COL[5355] = 1'b1;
assign COL[5356] = 1'b1;
assign COL[5357] = 1'b1;
assign COL[5358] = 1'b1;
assign COL[5359] = 1'b1;
assign COL[5360] = 1'b1;
assign COL[5361] = 1'b1;
assign COL[5362] = 1'b1;
assign COL[5363] = 1'b1;
assign COL[5364] = 1'b1;
assign COL[5365] = 1'b1;
assign COL[5366] = 1'b1;
assign COL[5367] = 1'b1;
assign COL[5368] = 1'b1;
assign COL[5369] = 1'b1;
assign COL[5370] = 1'b1;
assign COL[5371] = 1'b1;
assign COL[5372] = 1'b1;
assign COL[5373] = 1'b1;
assign COL[5374] = 1'b1;
assign COL[5375] = 1'b0;
assign COL[5376] = 1'b0;
assign COL[5377] = 1'b0;
assign COL[5378] = 1'b0;
assign COL[5379] = 1'b0;
assign COL[5380] = 1'b0;
assign COL[5381] = 1'b0;
assign COL[5382] = 1'b0;
assign COL[5383] = 1'b0;
assign COL[5384] = 1'b0;
assign COL[5385] = 1'b0;
assign COL[5386] = 1'b0;
assign COL[5387] = 1'b0;
assign COL[5388] = 1'b0;
assign COL[5389] = 1'b0;
assign COL[5390] = 1'b0;
assign COL[5391] = 1'b0;
assign COL[5392] = 1'b0;
assign COL[5393] = 1'b0;
assign COL[5394] = 1'b0;
assign COL[5395] = 1'b0;
assign COL[5396] = 1'b0;
assign COL[5397] = 1'b0;
assign COL[5398] = 1'b0;
assign COL[5399] = 1'b0;
assign COL[5400] = 1'b0;
assign COL[5401] = 1'b0;
assign COL[5402] = 1'b0;
assign COL[5403] = 1'b0;
assign COL[5404] = 1'b0;
assign COL[5405] = 1'b0;
assign COL[5406] = 1'b0;
assign COL[5407] = 1'b1;
assign COL[5408] = 1'b0;
assign COL[5409] = 1'b1;
assign COL[5410] = 1'b0;
assign COL[5411] = 1'b0;
assign COL[5412] = 1'b0;
assign COL[5413] = 1'b0;
assign COL[5414] = 1'b0;
assign COL[5415] = 1'b0;
assign COL[5416] = 1'b0;
assign COL[5417] = 1'b0;
assign COL[5418] = 1'b0;
assign COL[5419] = 1'b0;
assign COL[5420] = 1'b0;
assign COL[5421] = 1'b0;
assign COL[5422] = 1'b0;
assign COL[5423] = 1'b0;
assign COL[5424] = 1'b0;
assign COL[5425] = 1'b0;
assign COL[5426] = 1'b0;
assign COL[5427] = 1'b0;
assign COL[5428] = 1'b0;
assign COL[5429] = 1'b0;
assign COL[5430] = 1'b0;
assign COL[5431] = 1'b0;
assign COL[5432] = 1'b0;
assign COL[5433] = 1'b0;
assign COL[5434] = 1'b0;
assign COL[5435] = 1'b0;
assign COL[5436] = 1'b0;
assign COL[5437] = 1'b0;
assign COL[5438] = 1'b0;
assign COL[5439] = 1'b0;
assign COL[5440] = 1'b0;
assign COL[5441] = 1'b1;
assign COL[5442] = 1'b1;
assign COL[5443] = 1'b1;
assign COL[5444] = 1'b1;
assign COL[5445] = 1'b1;
assign COL[5446] = 1'b0;
assign COL[5447] = 1'b0;
assign COL[5448] = 1'b0;
assign COL[5449] = 1'b0;
assign COL[5450] = 1'b0;
assign COL[5451] = 1'b0;
assign COL[5452] = 1'b0;
assign COL[5453] = 1'b0;
assign COL[5454] = 1'b0;
assign COL[5455] = 1'b0;
assign COL[5456] = 1'b1;
assign COL[5457] = 1'b1;
assign COL[5458] = 1'b1;
assign COL[5459] = 1'b1;
assign COL[5460] = 1'b0;
assign COL[5461] = 1'b0;
assign COL[5462] = 1'b0;
assign COL[5463] = 1'b0;
assign COL[5464] = 1'b0;
assign COL[5465] = 1'b0;
assign COL[5466] = 1'b0;
assign COL[5467] = 1'b0;
assign COL[5468] = 1'b0;
assign COL[5469] = 1'b0;
assign COL[5470] = 1'b0;
assign COL[5471] = 1'b0;
assign COL[5472] = 1'b0;
assign COL[5473] = 1'b0;
assign COL[5474] = 1'b0;
assign COL[5475] = 1'b0;
assign COL[5476] = 1'b0;
assign COL[5477] = 1'b0;
assign COL[5478] = 1'b0;
assign COL[5479] = 1'b0;
assign COL[5480] = 1'b1;
assign COL[5481] = 1'b1;
assign COL[5482] = 1'b1;
assign COL[5483] = 1'b1;
assign COL[5484] = 1'b0;
assign COL[5485] = 1'b0;
assign COL[5486] = 1'b0;
assign COL[5487] = 1'b0;
assign COL[5488] = 1'b0;
assign COL[5489] = 1'b0;
assign COL[5490] = 1'b0;
assign COL[5491] = 1'b0;
assign COL[5492] = 1'b0;
assign COL[5493] = 1'b0;
assign COL[5494] = 1'b0;
assign COL[5495] = 1'b0;
assign COL[5496] = 1'b0;
assign COL[5497] = 1'b0;
assign COL[5498] = 1'b0;
assign COL[5499] = 1'b0;
assign COL[5500] = 1'b0;
assign COL[5501] = 1'b1;
assign COL[5502] = 1'b1;
assign COL[5503] = 1'b1;
assign COL[5504] = 1'b1;
assign COL[5505] = 1'b1;
assign COL[5506] = 1'b1;
assign COL[5507] = 1'b1;
assign COL[5508] = 1'b1;
assign COL[5509] = 1'b1;
assign COL[5510] = 1'b1;
assign COL[5511] = 1'b1;
assign COL[5512] = 1'b1;
assign COL[5513] = 1'b1;
assign COL[5514] = 1'b1;
assign COL[5515] = 1'b1;
assign COL[5516] = 1'b1;
assign COL[5517] = 1'b1;
assign COL[5518] = 1'b1;
assign COL[5519] = 1'b1;
assign COL[5520] = 1'b1;
assign COL[5521] = 1'b1;
assign COL[5522] = 1'b1;
assign COL[5523] = 1'b1;
assign COL[5524] = 1'b1;
assign COL[5525] = 1'b1;
assign COL[5526] = 1'b1;
assign COL[5527] = 1'b1;
assign COL[5528] = 1'b1;
assign COL[5529] = 1'b1;
assign COL[5530] = 1'b1;
assign COL[5531] = 1'b1;
assign COL[5532] = 1'b1;
assign COL[5533] = 1'b1;
assign COL[5534] = 1'b1;
assign COL[5535] = 1'b0;
assign COL[5536] = 1'b0;
assign COL[5537] = 1'b0;
assign COL[5538] = 1'b0;
assign COL[5539] = 1'b0;
assign COL[5540] = 1'b0;
assign COL[5541] = 1'b0;
assign COL[5542] = 1'b0;
assign COL[5543] = 1'b0;
assign COL[5544] = 1'b0;
assign COL[5545] = 1'b0;
assign COL[5546] = 1'b0;
assign COL[5547] = 1'b0;
assign COL[5548] = 1'b0;
assign COL[5549] = 1'b0;
assign COL[5550] = 1'b0;
assign COL[5551] = 1'b0;
assign COL[5552] = 1'b0;
assign COL[5553] = 1'b0;
assign COL[5554] = 1'b0;
assign COL[5555] = 1'b0;
assign COL[5556] = 1'b0;
assign COL[5557] = 1'b0;
assign COL[5558] = 1'b0;
assign COL[5559] = 1'b0;
assign COL[5560] = 1'b0;
assign COL[5561] = 1'b0;
assign COL[5562] = 1'b0;
assign COL[5563] = 1'b0;
assign COL[5564] = 1'b0;
assign COL[5565] = 1'b1;
assign COL[5566] = 1'b1;
assign COL[5567] = 1'b0;
assign COL[5568] = 1'b0;
assign COL[5569] = 1'b1;
assign COL[5570] = 1'b0;
assign COL[5571] = 1'b0;
assign COL[5572] = 1'b0;
assign COL[5573] = 1'b0;
assign COL[5574] = 1'b0;
assign COL[5575] = 1'b0;
assign COL[5576] = 1'b0;
assign COL[5577] = 1'b0;
assign COL[5578] = 1'b0;
assign COL[5579] = 1'b0;
assign COL[5580] = 1'b0;
assign COL[5581] = 1'b0;
assign COL[5582] = 1'b0;
assign COL[5583] = 1'b0;
assign COL[5584] = 1'b0;
assign COL[5585] = 1'b0;
assign COL[5586] = 1'b0;
assign COL[5587] = 1'b0;
assign COL[5588] = 1'b0;
assign COL[5589] = 1'b0;
assign COL[5590] = 1'b0;
assign COL[5591] = 1'b0;
assign COL[5592] = 1'b0;
assign COL[5593] = 1'b0;
assign COL[5594] = 1'b0;
assign COL[5595] = 1'b0;
assign COL[5596] = 1'b0;
assign COL[5597] = 1'b0;
assign COL[5598] = 1'b0;
assign COL[5599] = 1'b0;
assign COL[5600] = 1'b0;
assign COL[5601] = 1'b1;
assign COL[5602] = 1'b1;
assign COL[5603] = 1'b1;
assign COL[5604] = 1'b1;
assign COL[5605] = 1'b1;
assign COL[5606] = 1'b0;
assign COL[5607] = 1'b0;
assign COL[5608] = 1'b0;
assign COL[5609] = 1'b0;
assign COL[5610] = 1'b0;
assign COL[5611] = 1'b0;
assign COL[5612] = 1'b0;
assign COL[5613] = 1'b0;
assign COL[5614] = 1'b0;
assign COL[5615] = 1'b0;
assign COL[5616] = 1'b1;
assign COL[5617] = 1'b1;
assign COL[5618] = 1'b1;
assign COL[5619] = 1'b1;
assign COL[5620] = 1'b0;
assign COL[5621] = 1'b0;
assign COL[5622] = 1'b0;
assign COL[5623] = 1'b0;
assign COL[5624] = 1'b0;
assign COL[5625] = 1'b0;
assign COL[5626] = 1'b0;
assign COL[5627] = 1'b0;
assign COL[5628] = 1'b0;
assign COL[5629] = 1'b0;
assign COL[5630] = 1'b0;
assign COL[5631] = 1'b0;
assign COL[5632] = 1'b0;
assign COL[5633] = 1'b0;
assign COL[5634] = 1'b0;
assign COL[5635] = 1'b0;
assign COL[5636] = 1'b0;
assign COL[5637] = 1'b0;
assign COL[5638] = 1'b0;
assign COL[5639] = 1'b0;
assign COL[5640] = 1'b1;
assign COL[5641] = 1'b1;
assign COL[5642] = 1'b1;
assign COL[5643] = 1'b1;
assign COL[5644] = 1'b0;
assign COL[5645] = 1'b0;
assign COL[5646] = 1'b0;
assign COL[5647] = 1'b0;
assign COL[5648] = 1'b0;
assign COL[5649] = 1'b0;
assign COL[5650] = 1'b0;
assign COL[5651] = 1'b0;
assign COL[5652] = 1'b0;
assign COL[5653] = 1'b0;
assign COL[5654] = 1'b0;
assign COL[5655] = 1'b0;
assign COL[5656] = 1'b0;
assign COL[5657] = 1'b0;
assign COL[5658] = 1'b0;
assign COL[5659] = 1'b0;
assign COL[5660] = 1'b0;
assign COL[5661] = 1'b1;
assign COL[5662] = 1'b1;
assign COL[5663] = 1'b1;
assign COL[5664] = 1'b1;
assign COL[5665] = 1'b1;
assign COL[5666] = 1'b1;
assign COL[5667] = 1'b1;
assign COL[5668] = 1'b1;
assign COL[5669] = 1'b1;
assign COL[5670] = 1'b1;
assign COL[5671] = 1'b1;
assign COL[5672] = 1'b1;
assign COL[5673] = 1'b1;
assign COL[5674] = 1'b1;
assign COL[5675] = 1'b1;
assign COL[5676] = 1'b1;
assign COL[5677] = 1'b1;
assign COL[5678] = 1'b1;
assign COL[5679] = 1'b1;
assign COL[5680] = 1'b1;
assign COL[5681] = 1'b1;
assign COL[5682] = 1'b1;
assign COL[5683] = 1'b1;
assign COL[5684] = 1'b1;
assign COL[5685] = 1'b1;
assign COL[5686] = 1'b1;
assign COL[5687] = 1'b1;
assign COL[5688] = 1'b1;
assign COL[5689] = 1'b1;
assign COL[5690] = 1'b1;
assign COL[5691] = 1'b1;
assign COL[5692] = 1'b1;
assign COL[5693] = 1'b1;
assign COL[5694] = 1'b1;
assign COL[5695] = 1'b0;
assign COL[5696] = 1'b0;
assign COL[5697] = 1'b0;
assign COL[5698] = 1'b0;
assign COL[5699] = 1'b0;
assign COL[5700] = 1'b0;
assign COL[5701] = 1'b0;
assign COL[5702] = 1'b0;
assign COL[5703] = 1'b0;
assign COL[5704] = 1'b0;
assign COL[5705] = 1'b0;
assign COL[5706] = 1'b0;
assign COL[5707] = 1'b0;
assign COL[5708] = 1'b0;
assign COL[5709] = 1'b0;
assign COL[5710] = 1'b0;
assign COL[5711] = 1'b0;
assign COL[5712] = 1'b0;
assign COL[5713] = 1'b0;
assign COL[5714] = 1'b0;
assign COL[5715] = 1'b0;
assign COL[5716] = 1'b0;
assign COL[5717] = 1'b0;
assign COL[5718] = 1'b0;
assign COL[5719] = 1'b0;
assign COL[5720] = 1'b0;
assign COL[5721] = 1'b0;
assign COL[5722] = 1'b0;
assign COL[5723] = 1'b0;
assign COL[5724] = 1'b0;
assign COL[5725] = 1'b0;
assign COL[5726] = 1'b0;
assign COL[5727] = 1'b0;
assign COL[5728] = 1'b0;
assign COL[5729] = 1'b0;
assign COL[5730] = 1'b0;
assign COL[5731] = 1'b0;
assign COL[5732] = 1'b0;
assign COL[5733] = 1'b0;
assign COL[5734] = 1'b0;
assign COL[5735] = 1'b0;
assign COL[5736] = 1'b0;
assign COL[5737] = 1'b0;
assign COL[5738] = 1'b0;
assign COL[5739] = 1'b0;
assign COL[5740] = 1'b0;
assign COL[5741] = 1'b0;
assign COL[5742] = 1'b0;
assign COL[5743] = 1'b0;
assign COL[5744] = 1'b0;
assign COL[5745] = 1'b0;
assign COL[5746] = 1'b0;
assign COL[5747] = 1'b0;
assign COL[5748] = 1'b0;
assign COL[5749] = 1'b0;
assign COL[5750] = 1'b0;
assign COL[5751] = 1'b0;
assign COL[5752] = 1'b0;
assign COL[5753] = 1'b0;
assign COL[5754] = 1'b0;
assign COL[5755] = 1'b0;
assign COL[5756] = 1'b0;
assign COL[5757] = 1'b0;
assign COL[5758] = 1'b0;
assign COL[5759] = 1'b0;
assign COL[5760] = 1'b0;
assign COL[5761] = 1'b1;
assign COL[5762] = 1'b1;
assign COL[5763] = 1'b1;
assign COL[5764] = 1'b1;
assign COL[5765] = 1'b1;
assign COL[5766] = 1'b0;
assign COL[5767] = 1'b0;
assign COL[5768] = 1'b0;
assign COL[5769] = 1'b0;
assign COL[5770] = 1'b0;
assign COL[5771] = 1'b0;
assign COL[5772] = 1'b0;
assign COL[5773] = 1'b0;
assign COL[5774] = 1'b0;
assign COL[5775] = 1'b0;
assign COL[5776] = 1'b1;
assign COL[5777] = 1'b1;
assign COL[5778] = 1'b1;
assign COL[5779] = 1'b1;
assign COL[5780] = 1'b0;
assign COL[5781] = 1'b0;
assign COL[5782] = 1'b0;
assign COL[5783] = 1'b0;
assign COL[5784] = 1'b0;
assign COL[5785] = 1'b0;
assign COL[5786] = 1'b0;
assign COL[5787] = 1'b0;
assign COL[5788] = 1'b0;
assign COL[5789] = 1'b0;
assign COL[5790] = 1'b0;
assign COL[5791] = 1'b0;
assign COL[5792] = 1'b0;
assign COL[5793] = 1'b0;
assign COL[5794] = 1'b0;
assign COL[5795] = 1'b0;
assign COL[5796] = 1'b0;
assign COL[5797] = 1'b0;
assign COL[5798] = 1'b0;
assign COL[5799] = 1'b0;
assign COL[5800] = 1'b1;
assign COL[5801] = 1'b1;
assign COL[5802] = 1'b1;
assign COL[5803] = 1'b1;
assign COL[5804] = 1'b0;
assign COL[5805] = 1'b0;
assign COL[5806] = 1'b0;
assign COL[5807] = 1'b0;
assign COL[5808] = 1'b0;
assign COL[5809] = 1'b0;
assign COL[5810] = 1'b0;
assign COL[5811] = 1'b0;
assign COL[5812] = 1'b0;
assign COL[5813] = 1'b0;
assign COL[5814] = 1'b0;
assign COL[5815] = 1'b0;
assign COL[5816] = 1'b0;
assign COL[5817] = 1'b0;
assign COL[5818] = 1'b0;
assign COL[5819] = 1'b0;
assign COL[5820] = 1'b0;
assign COL[5821] = 1'b1;
assign COL[5822] = 1'b1;
assign COL[5823] = 1'b1;
assign COL[5824] = 1'b1;
assign COL[5825] = 1'b1;
assign COL[5826] = 1'b1;
assign COL[5827] = 1'b1;
assign COL[5828] = 1'b1;
assign COL[5829] = 1'b1;
assign COL[5830] = 1'b1;
assign COL[5831] = 1'b1;
assign COL[5832] = 1'b1;
assign COL[5833] = 1'b1;
assign COL[5834] = 1'b1;
assign COL[5835] = 1'b1;
assign COL[5836] = 1'b1;
assign COL[5837] = 1'b1;
assign COL[5838] = 1'b1;
assign COL[5839] = 1'b1;
assign COL[5840] = 1'b1;
assign COL[5841] = 1'b1;
assign COL[5842] = 1'b1;
assign COL[5843] = 1'b1;
assign COL[5844] = 1'b1;
assign COL[5845] = 1'b1;
assign COL[5846] = 1'b1;
assign COL[5847] = 1'b1;
assign COL[5848] = 1'b1;
assign COL[5849] = 1'b1;
assign COL[5850] = 1'b1;
assign COL[5851] = 1'b1;
assign COL[5852] = 1'b1;
assign COL[5853] = 1'b1;
assign COL[5854] = 1'b1;
assign COL[5855] = 1'b0;
assign COL[5856] = 1'b0;
assign COL[5857] = 1'b0;
assign COL[5858] = 1'b0;
assign COL[5859] = 1'b0;
assign COL[5860] = 1'b0;
assign COL[5861] = 1'b0;
assign COL[5862] = 1'b0;
assign COL[5863] = 1'b0;
assign COL[5864] = 1'b0;
assign COL[5865] = 1'b0;
assign COL[5866] = 1'b0;
assign COL[5867] = 1'b0;
assign COL[5868] = 1'b0;
assign COL[5869] = 1'b0;
assign COL[5870] = 1'b0;
assign COL[5871] = 1'b0;
assign COL[5872] = 1'b0;
assign COL[5873] = 1'b0;
assign COL[5874] = 1'b0;
assign COL[5875] = 1'b0;
assign COL[5876] = 1'b0;
assign COL[5877] = 1'b0;
assign COL[5878] = 1'b0;
assign COL[5879] = 1'b0;
assign COL[5880] = 1'b0;
assign COL[5881] = 1'b0;
assign COL[5882] = 1'b0;
assign COL[5883] = 1'b0;
assign COL[5884] = 1'b0;
assign COL[5885] = 1'b0;
assign COL[5886] = 1'b0;
assign COL[5887] = 1'b1;
assign COL[5888] = 1'b0;
assign COL[5889] = 1'b0;
assign COL[5890] = 1'b0;
assign COL[5891] = 1'b0;
assign COL[5892] = 1'b0;
assign COL[5893] = 1'b0;
assign COL[5894] = 1'b0;
assign COL[5895] = 1'b0;
assign COL[5896] = 1'b0;
assign COL[5897] = 1'b0;
assign COL[5898] = 1'b0;
assign COL[5899] = 1'b0;
assign COL[5900] = 1'b0;
assign COL[5901] = 1'b0;
assign COL[5902] = 1'b0;
assign COL[5903] = 1'b0;
assign COL[5904] = 1'b0;
assign COL[5905] = 1'b0;
assign COL[5906] = 1'b0;
assign COL[5907] = 1'b0;
assign COL[5908] = 1'b0;
assign COL[5909] = 1'b0;
assign COL[5910] = 1'b0;
assign COL[5911] = 1'b0;
assign COL[5912] = 1'b0;
assign COL[5913] = 1'b0;
assign COL[5914] = 1'b0;
assign COL[5915] = 1'b0;
assign COL[5916] = 1'b0;
assign COL[5917] = 1'b0;
assign COL[5918] = 1'b0;
assign COL[5919] = 1'b0;
assign COL[5920] = 1'b0;
assign COL[5921] = 1'b1;
assign COL[5922] = 1'b1;
assign COL[5923] = 1'b1;
assign COL[5924] = 1'b1;
assign COL[5925] = 1'b1;
assign COL[5926] = 1'b0;
assign COL[5927] = 1'b0;
assign COL[5928] = 1'b0;
assign COL[5929] = 1'b0;
assign COL[5930] = 1'b0;
assign COL[5931] = 1'b0;
assign COL[5932] = 1'b0;
assign COL[5933] = 1'b0;
assign COL[5934] = 1'b0;
assign COL[5935] = 1'b0;
assign COL[5936] = 1'b1;
assign COL[5937] = 1'b1;
assign COL[5938] = 1'b1;
assign COL[5939] = 1'b1;
assign COL[5940] = 1'b0;
assign COL[5941] = 1'b0;
assign COL[5942] = 1'b0;
assign COL[5943] = 1'b0;
assign COL[5944] = 1'b0;
assign COL[5945] = 1'b0;
assign COL[5946] = 1'b0;
assign COL[5947] = 1'b0;
assign COL[5948] = 1'b0;
assign COL[5949] = 1'b0;
assign COL[5950] = 1'b0;
assign COL[5951] = 1'b0;
assign COL[5952] = 1'b0;
assign COL[5953] = 1'b0;
assign COL[5954] = 1'b0;
assign COL[5955] = 1'b0;
assign COL[5956] = 1'b0;
assign COL[5957] = 1'b0;
assign COL[5958] = 1'b0;
assign COL[5959] = 1'b0;
assign COL[5960] = 1'b1;
assign COL[5961] = 1'b1;
assign COL[5962] = 1'b1;
assign COL[5963] = 1'b1;
assign COL[5964] = 1'b0;
assign COL[5965] = 1'b0;
assign COL[5966] = 1'b0;
assign COL[5967] = 1'b0;
assign COL[5968] = 1'b0;
assign COL[5969] = 1'b0;
assign COL[5970] = 1'b0;
assign COL[5971] = 1'b0;
assign COL[5972] = 1'b0;
assign COL[5973] = 1'b0;
assign COL[5974] = 1'b0;
assign COL[5975] = 1'b0;
assign COL[5976] = 1'b0;
assign COL[5977] = 1'b0;
assign COL[5978] = 1'b0;
assign COL[5979] = 1'b0;
assign COL[5980] = 1'b0;
assign COL[5981] = 1'b1;
assign COL[5982] = 1'b1;
assign COL[5983] = 1'b1;
assign COL[5984] = 1'b1;
assign COL[5985] = 1'b1;
assign COL[5986] = 1'b1;
assign COL[5987] = 1'b1;
assign COL[5988] = 1'b1;
assign COL[5989] = 1'b1;
assign COL[5990] = 1'b1;
assign COL[5991] = 1'b1;
assign COL[5992] = 1'b1;
assign COL[5993] = 1'b1;
assign COL[5994] = 1'b1;
assign COL[5995] = 1'b1;
assign COL[5996] = 1'b1;
assign COL[5997] = 1'b1;
assign COL[5998] = 1'b1;
assign COL[5999] = 1'b1;
assign COL[6000] = 1'b1;
assign COL[6001] = 1'b1;
assign COL[6002] = 1'b1;
assign COL[6003] = 1'b1;
assign COL[6004] = 1'b1;
assign COL[6005] = 1'b1;
assign COL[6006] = 1'b1;
assign COL[6007] = 1'b1;
assign COL[6008] = 1'b1;
assign COL[6009] = 1'b1;
assign COL[6010] = 1'b1;
assign COL[6011] = 1'b1;
assign COL[6012] = 1'b1;
assign COL[6013] = 1'b1;
assign COL[6014] = 1'b1;
assign COL[6015] = 1'b0;
assign COL[6016] = 1'b0;
assign COL[6017] = 1'b0;
assign COL[6018] = 1'b0;
assign COL[6019] = 1'b0;
assign COL[6020] = 1'b0;
assign COL[6021] = 1'b0;
assign COL[6022] = 1'b0;
assign COL[6023] = 1'b0;
assign COL[6024] = 1'b0;
assign COL[6025] = 1'b0;
assign COL[6026] = 1'b0;
assign COL[6027] = 1'b0;
assign COL[6028] = 1'b0;
assign COL[6029] = 1'b0;
assign COL[6030] = 1'b0;
assign COL[6031] = 1'b0;
assign COL[6032] = 1'b0;
assign COL[6033] = 1'b0;
assign COL[6034] = 1'b0;
assign COL[6035] = 1'b0;
assign COL[6036] = 1'b0;
assign COL[6037] = 1'b0;
assign COL[6038] = 1'b0;
assign COL[6039] = 1'b0;
assign COL[6040] = 1'b0;
assign COL[6041] = 1'b0;
assign COL[6042] = 1'b0;
assign COL[6043] = 1'b0;
assign COL[6044] = 1'b0;
assign COL[6045] = 1'b0;
assign COL[6046] = 1'b0;
assign COL[6047] = 1'b0;
assign COL[6048] = 1'b0;
assign COL[6049] = 1'b0;
assign COL[6050] = 1'b0;
assign COL[6051] = 1'b0;
assign COL[6052] = 1'b0;
assign COL[6053] = 1'b0;
assign COL[6054] = 1'b0;
assign COL[6055] = 1'b0;
assign COL[6056] = 1'b0;
assign COL[6057] = 1'b0;
assign COL[6058] = 1'b0;
assign COL[6059] = 1'b0;
assign COL[6060] = 1'b0;
assign COL[6061] = 1'b0;
assign COL[6062] = 1'b0;
assign COL[6063] = 1'b0;
assign COL[6064] = 1'b0;
assign COL[6065] = 1'b0;
assign COL[6066] = 1'b0;
assign COL[6067] = 1'b0;
assign COL[6068] = 1'b0;
assign COL[6069] = 1'b0;
assign COL[6070] = 1'b0;
assign COL[6071] = 1'b0;
assign COL[6072] = 1'b0;
assign COL[6073] = 1'b0;
assign COL[6074] = 1'b0;
assign COL[6075] = 1'b0;
assign COL[6076] = 1'b0;
assign COL[6077] = 1'b0;
assign COL[6078] = 1'b0;
assign COL[6079] = 1'b0;
assign COL[6080] = 1'b0;
assign COL[6081] = 1'b1;
assign COL[6082] = 1'b1;
assign COL[6083] = 1'b1;
assign COL[6084] = 1'b1;
assign COL[6085] = 1'b1;
assign COL[6086] = 1'b0;
assign COL[6087] = 1'b0;
assign COL[6088] = 1'b0;
assign COL[6089] = 1'b0;
assign COL[6090] = 1'b0;
assign COL[6091] = 1'b0;
assign COL[6092] = 1'b0;
assign COL[6093] = 1'b0;
assign COL[6094] = 1'b0;
assign COL[6095] = 1'b0;
assign COL[6096] = 1'b1;
assign COL[6097] = 1'b1;
assign COL[6098] = 1'b1;
assign COL[6099] = 1'b1;
assign COL[6100] = 1'b0;
assign COL[6101] = 1'b0;
assign COL[6102] = 1'b0;
assign COL[6103] = 1'b0;
assign COL[6104] = 1'b0;
assign COL[6105] = 1'b0;
assign COL[6106] = 1'b0;
assign COL[6107] = 1'b0;
assign COL[6108] = 1'b0;
assign COL[6109] = 1'b0;
assign COL[6110] = 1'b0;
assign COL[6111] = 1'b0;
assign COL[6112] = 1'b0;
assign COL[6113] = 1'b0;
assign COL[6114] = 1'b0;
assign COL[6115] = 1'b0;
assign COL[6116] = 1'b0;
assign COL[6117] = 1'b0;
assign COL[6118] = 1'b0;
assign COL[6119] = 1'b0;
assign COL[6120] = 1'b1;
assign COL[6121] = 1'b1;
assign COL[6122] = 1'b1;
assign COL[6123] = 1'b1;
assign COL[6124] = 1'b0;
assign COL[6125] = 1'b0;
assign COL[6126] = 1'b0;
assign COL[6127] = 1'b0;
assign COL[6128] = 1'b0;
assign COL[6129] = 1'b0;
assign COL[6130] = 1'b0;
assign COL[6131] = 1'b0;
assign COL[6132] = 1'b0;
assign COL[6133] = 1'b0;
assign COL[6134] = 1'b0;
assign COL[6135] = 1'b0;
assign COL[6136] = 1'b0;
assign COL[6137] = 1'b0;
assign COL[6138] = 1'b0;
assign COL[6139] = 1'b0;
assign COL[6140] = 1'b0;
assign COL[6141] = 1'b0;
assign COL[6142] = 1'b0;
assign COL[6143] = 1'b0;
assign COL[6144] = 1'b0;
assign COL[6145] = 1'b0;
assign COL[6146] = 1'b0;
assign COL[6147] = 1'b0;
assign COL[6148] = 1'b0;
assign COL[6149] = 1'b0;
assign COL[6150] = 1'b0;
assign COL[6151] = 1'b0;
assign COL[6152] = 1'b0;
assign COL[6153] = 1'b0;
assign COL[6154] = 1'b0;
assign COL[6155] = 1'b0;
assign COL[6156] = 1'b0;
assign COL[6157] = 1'b0;
assign COL[6158] = 1'b0;
assign COL[6159] = 1'b0;
assign COL[6160] = 1'b0;
assign COL[6161] = 1'b0;
assign COL[6162] = 1'b0;
assign COL[6163] = 1'b0;
assign COL[6164] = 1'b0;
assign COL[6165] = 1'b0;
assign COL[6166] = 1'b0;
assign COL[6167] = 1'b0;
assign COL[6168] = 1'b0;
assign COL[6169] = 1'b0;
assign COL[6170] = 1'b1;
assign COL[6171] = 1'b1;
assign COL[6172] = 1'b1;
assign COL[6173] = 1'b1;
assign COL[6174] = 1'b1;
assign COL[6175] = 1'b0;
assign COL[6176] = 1'b0;
assign COL[6177] = 1'b0;
assign COL[6178] = 1'b0;
assign COL[6179] = 1'b0;
assign COL[6180] = 1'b0;
assign COL[6181] = 1'b0;
assign COL[6182] = 1'b0;
assign COL[6183] = 1'b0;
assign COL[6184] = 1'b0;
assign COL[6185] = 1'b0;
assign COL[6186] = 1'b0;
assign COL[6187] = 1'b0;
assign COL[6188] = 1'b0;
assign COL[6189] = 1'b0;
assign COL[6190] = 1'b0;
assign COL[6191] = 1'b0;
assign COL[6192] = 1'b0;
assign COL[6193] = 1'b0;
assign COL[6194] = 1'b0;
assign COL[6195] = 1'b0;
assign COL[6196] = 1'b0;
assign COL[6197] = 1'b0;
assign COL[6198] = 1'b0;
assign COL[6199] = 1'b0;
assign COL[6200] = 1'b0;
assign COL[6201] = 1'b0;
assign COL[6202] = 1'b0;
assign COL[6203] = 1'b0;
assign COL[6204] = 1'b0;
assign COL[6205] = 1'b0;
assign COL[6206] = 1'b0;
assign COL[6207] = 1'b0;
assign COL[6208] = 1'b0;
assign COL[6209] = 1'b0;
assign COL[6210] = 1'b0;
assign COL[6211] = 1'b0;
assign COL[6212] = 1'b0;
assign COL[6213] = 1'b0;
assign COL[6214] = 1'b0;
assign COL[6215] = 1'b0;
assign COL[6216] = 1'b0;
assign COL[6217] = 1'b0;
assign COL[6218] = 1'b0;
assign COL[6219] = 1'b0;
assign COL[6220] = 1'b0;
assign COL[6221] = 1'b0;
assign COL[6222] = 1'b0;
assign COL[6223] = 1'b0;
assign COL[6224] = 1'b0;
assign COL[6225] = 1'b0;
assign COL[6226] = 1'b0;
assign COL[6227] = 1'b0;
assign COL[6228] = 1'b0;
assign COL[6229] = 1'b0;
assign COL[6230] = 1'b0;
assign COL[6231] = 1'b0;
assign COL[6232] = 1'b0;
assign COL[6233] = 1'b0;
assign COL[6234] = 1'b0;
assign COL[6235] = 1'b0;
assign COL[6236] = 1'b0;
assign COL[6237] = 1'b0;
assign COL[6238] = 1'b0;
assign COL[6239] = 1'b0;
assign COL[6240] = 1'b0;
assign COL[6241] = 1'b1;
assign COL[6242] = 1'b1;
assign COL[6243] = 1'b1;
assign COL[6244] = 1'b1;
assign COL[6245] = 1'b1;
assign COL[6246] = 1'b0;
assign COL[6247] = 1'b0;
assign COL[6248] = 1'b0;
assign COL[6249] = 1'b0;
assign COL[6250] = 1'b0;
assign COL[6251] = 1'b0;
assign COL[6252] = 1'b0;
assign COL[6253] = 1'b0;
assign COL[6254] = 1'b0;
assign COL[6255] = 1'b0;
assign COL[6256] = 1'b1;
assign COL[6257] = 1'b1;
assign COL[6258] = 1'b1;
assign COL[6259] = 1'b1;
assign COL[6260] = 1'b0;
assign COL[6261] = 1'b0;
assign COL[6262] = 1'b0;
assign COL[6263] = 1'b0;
assign COL[6264] = 1'b0;
assign COL[6265] = 1'b0;
assign COL[6266] = 1'b0;
assign COL[6267] = 1'b0;
assign COL[6268] = 1'b0;
assign COL[6269] = 1'b0;
assign COL[6270] = 1'b0;
assign COL[6271] = 1'b0;
assign COL[6272] = 1'b0;
assign COL[6273] = 1'b0;
assign COL[6274] = 1'b0;
assign COL[6275] = 1'b0;
assign COL[6276] = 1'b0;
assign COL[6277] = 1'b0;
assign COL[6278] = 1'b0;
assign COL[6279] = 1'b0;
assign COL[6280] = 1'b1;
assign COL[6281] = 1'b1;
assign COL[6282] = 1'b1;
assign COL[6283] = 1'b1;
assign COL[6284] = 1'b0;
assign COL[6285] = 1'b0;
assign COL[6286] = 1'b0;
assign COL[6287] = 1'b0;
assign COL[6288] = 1'b0;
assign COL[6289] = 1'b0;
assign COL[6290] = 1'b0;
assign COL[6291] = 1'b0;
assign COL[6292] = 1'b0;
assign COL[6293] = 1'b0;
assign COL[6294] = 1'b0;
assign COL[6295] = 1'b0;
assign COL[6296] = 1'b0;
assign COL[6297] = 1'b0;
assign COL[6298] = 1'b0;
assign COL[6299] = 1'b0;
assign COL[6300] = 1'b0;
assign COL[6301] = 1'b0;
assign COL[6302] = 1'b0;
assign COL[6303] = 1'b0;
assign COL[6304] = 1'b0;
assign COL[6305] = 1'b0;
assign COL[6306] = 1'b0;
assign COL[6307] = 1'b0;
assign COL[6308] = 1'b0;
assign COL[6309] = 1'b0;
assign COL[6310] = 1'b0;
assign COL[6311] = 1'b0;
assign COL[6312] = 1'b0;
assign COL[6313] = 1'b0;
assign COL[6314] = 1'b0;
assign COL[6315] = 1'b0;
assign COL[6316] = 1'b0;
assign COL[6317] = 1'b0;
assign COL[6318] = 1'b0;
assign COL[6319] = 1'b0;
assign COL[6320] = 1'b0;
assign COL[6321] = 1'b0;
assign COL[6322] = 1'b0;
assign COL[6323] = 1'b0;
assign COL[6324] = 1'b0;
assign COL[6325] = 1'b0;
assign COL[6326] = 1'b0;
assign COL[6327] = 1'b0;
assign COL[6328] = 1'b0;
assign COL[6329] = 1'b0;
assign COL[6330] = 1'b1;
assign COL[6331] = 1'b1;
assign COL[6332] = 1'b1;
assign COL[6333] = 1'b1;
assign COL[6334] = 1'b1;
assign COL[6335] = 1'b0;
assign COL[6336] = 1'b0;
assign COL[6337] = 1'b0;
assign COL[6338] = 1'b0;
assign COL[6339] = 1'b0;
assign COL[6340] = 1'b0;
assign COL[6341] = 1'b0;
assign COL[6342] = 1'b0;
assign COL[6343] = 1'b0;
assign COL[6344] = 1'b0;
assign COL[6345] = 1'b0;
assign COL[6346] = 1'b0;
assign COL[6347] = 1'b0;
assign COL[6348] = 1'b0;
assign COL[6349] = 1'b0;
assign COL[6350] = 1'b0;
assign COL[6351] = 1'b0;
assign COL[6352] = 1'b0;
assign COL[6353] = 1'b0;
assign COL[6354] = 1'b0;
assign COL[6355] = 1'b0;
assign COL[6356] = 1'b0;
assign COL[6357] = 1'b0;
assign COL[6358] = 1'b0;
assign COL[6359] = 1'b0;
assign COL[6360] = 1'b0;
assign COL[6361] = 1'b0;
assign COL[6362] = 1'b0;
assign COL[6363] = 1'b0;
assign COL[6364] = 1'b0;
assign COL[6365] = 1'b0;
assign COL[6366] = 1'b0;
assign COL[6367] = 1'b0;
assign COL[6368] = 1'b0;
assign COL[6369] = 1'b0;
assign COL[6370] = 1'b0;
assign COL[6371] = 1'b0;
assign COL[6372] = 1'b0;
assign COL[6373] = 1'b0;
assign COL[6374] = 1'b0;
assign COL[6375] = 1'b0;
assign COL[6376] = 1'b0;
assign COL[6377] = 1'b0;
assign COL[6378] = 1'b0;
assign COL[6379] = 1'b0;
assign COL[6380] = 1'b0;
assign COL[6381] = 1'b0;
assign COL[6382] = 1'b0;
assign COL[6383] = 1'b0;
assign COL[6384] = 1'b0;
assign COL[6385] = 1'b0;
assign COL[6386] = 1'b0;
assign COL[6387] = 1'b0;
assign COL[6388] = 1'b0;
assign COL[6389] = 1'b0;
assign COL[6390] = 1'b0;
assign COL[6391] = 1'b0;
assign COL[6392] = 1'b0;
assign COL[6393] = 1'b0;
assign COL[6394] = 1'b0;
assign COL[6395] = 1'b0;
assign COL[6396] = 1'b0;
assign COL[6397] = 1'b0;
assign COL[6398] = 1'b0;
assign COL[6399] = 1'b0;
assign COL[6400] = 1'b0;
assign COL[6401] = 1'b1;
assign COL[6402] = 1'b1;
assign COL[6403] = 1'b1;
assign COL[6404] = 1'b1;
assign COL[6405] = 1'b1;
assign COL[6406] = 1'b0;
assign COL[6407] = 1'b0;
assign COL[6408] = 1'b0;
assign COL[6409] = 1'b0;
assign COL[6410] = 1'b0;
assign COL[6411] = 1'b0;
assign COL[6412] = 1'b0;
assign COL[6413] = 1'b0;
assign COL[6414] = 1'b0;
assign COL[6415] = 1'b0;
assign COL[6416] = 1'b1;
assign COL[6417] = 1'b1;
assign COL[6418] = 1'b1;
assign COL[6419] = 1'b1;
assign COL[6420] = 1'b0;
assign COL[6421] = 1'b0;
assign COL[6422] = 1'b0;
assign COL[6423] = 1'b0;
assign COL[6424] = 1'b0;
assign COL[6425] = 1'b0;
assign COL[6426] = 1'b0;
assign COL[6427] = 1'b0;
assign COL[6428] = 1'b0;
assign COL[6429] = 1'b0;
assign COL[6430] = 1'b0;
assign COL[6431] = 1'b0;
assign COL[6432] = 1'b0;
assign COL[6433] = 1'b0;
assign COL[6434] = 1'b0;
assign COL[6435] = 1'b0;
assign COL[6436] = 1'b0;
assign COL[6437] = 1'b0;
assign COL[6438] = 1'b0;
assign COL[6439] = 1'b0;
assign COL[6440] = 1'b1;
assign COL[6441] = 1'b1;
assign COL[6442] = 1'b1;
assign COL[6443] = 1'b1;
assign COL[6444] = 1'b0;
assign COL[6445] = 1'b0;
assign COL[6446] = 1'b0;
assign COL[6447] = 1'b0;
assign COL[6448] = 1'b0;
assign COL[6449] = 1'b0;
assign COL[6450] = 1'b0;
assign COL[6451] = 1'b0;
assign COL[6452] = 1'b0;
assign COL[6453] = 1'b0;
assign COL[6454] = 1'b0;
assign COL[6455] = 1'b0;
assign COL[6456] = 1'b0;
assign COL[6457] = 1'b0;
assign COL[6458] = 1'b0;
assign COL[6459] = 1'b0;
assign COL[6460] = 1'b0;
assign COL[6461] = 1'b0;
assign COL[6462] = 1'b0;
assign COL[6463] = 1'b0;
assign COL[6464] = 1'b0;
assign COL[6465] = 1'b0;
assign COL[6466] = 1'b0;
assign COL[6467] = 1'b0;
assign COL[6468] = 1'b0;
assign COL[6469] = 1'b0;
assign COL[6470] = 1'b0;
assign COL[6471] = 1'b0;
assign COL[6472] = 1'b0;
assign COL[6473] = 1'b0;
assign COL[6474] = 1'b0;
assign COL[6475] = 1'b0;
assign COL[6476] = 1'b0;
assign COL[6477] = 1'b0;
assign COL[6478] = 1'b0;
assign COL[6479] = 1'b0;
assign COL[6480] = 1'b0;
assign COL[6481] = 1'b0;
assign COL[6482] = 1'b0;
assign COL[6483] = 1'b0;
assign COL[6484] = 1'b0;
assign COL[6485] = 1'b0;
assign COL[6486] = 1'b0;
assign COL[6487] = 1'b0;
assign COL[6488] = 1'b0;
assign COL[6489] = 1'b0;
assign COL[6490] = 1'b1;
assign COL[6491] = 1'b1;
assign COL[6492] = 1'b1;
assign COL[6493] = 1'b1;
assign COL[6494] = 1'b1;
assign COL[6495] = 1'b0;
assign COL[6496] = 1'b0;
assign COL[6497] = 1'b0;
assign COL[6498] = 1'b0;
assign COL[6499] = 1'b0;
assign COL[6500] = 1'b0;
assign COL[6501] = 1'b0;
assign COL[6502] = 1'b0;
assign COL[6503] = 1'b0;
assign COL[6504] = 1'b0;
assign COL[6505] = 1'b0;
assign COL[6506] = 1'b0;
assign COL[6507] = 1'b0;
assign COL[6508] = 1'b0;
assign COL[6509] = 1'b0;
assign COL[6510] = 1'b0;
assign COL[6511] = 1'b0;
assign COL[6512] = 1'b0;
assign COL[6513] = 1'b0;
assign COL[6514] = 1'b0;
assign COL[6515] = 1'b0;
assign COL[6516] = 1'b0;
assign COL[6517] = 1'b0;
assign COL[6518] = 1'b0;
assign COL[6519] = 1'b0;
assign COL[6520] = 1'b0;
assign COL[6521] = 1'b0;
assign COL[6522] = 1'b0;
assign COL[6523] = 1'b0;
assign COL[6524] = 1'b0;
assign COL[6525] = 1'b0;
assign COL[6526] = 1'b0;
assign COL[6527] = 1'b0;
assign COL[6528] = 1'b0;
assign COL[6529] = 1'b0;
assign COL[6530] = 1'b0;
assign COL[6531] = 1'b0;
assign COL[6532] = 1'b0;
assign COL[6533] = 1'b0;
assign COL[6534] = 1'b0;
assign COL[6535] = 1'b0;
assign COL[6536] = 1'b0;
assign COL[6537] = 1'b0;
assign COL[6538] = 1'b0;
assign COL[6539] = 1'b0;
assign COL[6540] = 1'b0;
assign COL[6541] = 1'b0;
assign COL[6542] = 1'b0;
assign COL[6543] = 1'b0;
assign COL[6544] = 1'b0;
assign COL[6545] = 1'b0;
assign COL[6546] = 1'b0;
assign COL[6547] = 1'b0;
assign COL[6548] = 1'b0;
assign COL[6549] = 1'b0;
assign COL[6550] = 1'b0;
assign COL[6551] = 1'b0;
assign COL[6552] = 1'b0;
assign COL[6553] = 1'b0;
assign COL[6554] = 1'b0;
assign COL[6555] = 1'b0;
assign COL[6556] = 1'b0;
assign COL[6557] = 1'b0;
assign COL[6558] = 1'b0;
assign COL[6559] = 1'b0;
assign COL[6560] = 1'b0;
assign COL[6561] = 1'b1;
assign COL[6562] = 1'b1;
assign COL[6563] = 1'b1;
assign COL[6564] = 1'b1;
assign COL[6565] = 1'b1;
assign COL[6566] = 1'b0;
assign COL[6567] = 1'b0;
assign COL[6568] = 1'b0;
assign COL[6569] = 1'b0;
assign COL[6570] = 1'b0;
assign COL[6571] = 1'b0;
assign COL[6572] = 1'b0;
assign COL[6573] = 1'b0;
assign COL[6574] = 1'b0;
assign COL[6575] = 1'b0;
assign COL[6576] = 1'b1;
assign COL[6577] = 1'b1;
assign COL[6578] = 1'b1;
assign COL[6579] = 1'b1;
assign COL[6580] = 1'b0;
assign COL[6581] = 1'b0;
assign COL[6582] = 1'b0;
assign COL[6583] = 1'b0;
assign COL[6584] = 1'b0;
assign COL[6585] = 1'b0;
assign COL[6586] = 1'b0;
assign COL[6587] = 1'b0;
assign COL[6588] = 1'b0;
assign COL[6589] = 1'b0;
assign COL[6590] = 1'b0;
assign COL[6591] = 1'b0;
assign COL[6592] = 1'b0;
assign COL[6593] = 1'b0;
assign COL[6594] = 1'b0;
assign COL[6595] = 1'b0;
assign COL[6596] = 1'b0;
assign COL[6597] = 1'b0;
assign COL[6598] = 1'b0;
assign COL[6599] = 1'b0;
assign COL[6600] = 1'b1;
assign COL[6601] = 1'b1;
assign COL[6602] = 1'b1;
assign COL[6603] = 1'b1;
assign COL[6604] = 1'b0;
assign COL[6605] = 1'b0;
assign COL[6606] = 1'b0;
assign COL[6607] = 1'b0;
assign COL[6608] = 1'b0;
assign COL[6609] = 1'b0;
assign COL[6610] = 1'b0;
assign COL[6611] = 1'b0;
assign COL[6612] = 1'b0;
assign COL[6613] = 1'b0;
assign COL[6614] = 1'b0;
assign COL[6615] = 1'b0;
assign COL[6616] = 1'b0;
assign COL[6617] = 1'b0;
assign COL[6618] = 1'b0;
assign COL[6619] = 1'b0;
assign COL[6620] = 1'b0;
assign COL[6621] = 1'b0;
assign COL[6622] = 1'b0;
assign COL[6623] = 1'b0;
assign COL[6624] = 1'b0;
assign COL[6625] = 1'b0;
assign COL[6626] = 1'b0;
assign COL[6627] = 1'b0;
assign COL[6628] = 1'b0;
assign COL[6629] = 1'b0;
assign COL[6630] = 1'b0;
assign COL[6631] = 1'b0;
assign COL[6632] = 1'b0;
assign COL[6633] = 1'b0;
assign COL[6634] = 1'b0;
assign COL[6635] = 1'b0;
assign COL[6636] = 1'b0;
assign COL[6637] = 1'b0;
assign COL[6638] = 1'b0;
assign COL[6639] = 1'b0;
assign COL[6640] = 1'b0;
assign COL[6641] = 1'b0;
assign COL[6642] = 1'b0;
assign COL[6643] = 1'b0;
assign COL[6644] = 1'b0;
assign COL[6645] = 1'b0;
assign COL[6646] = 1'b0;
assign COL[6647] = 1'b0;
assign COL[6648] = 1'b0;
assign COL[6649] = 1'b0;
assign COL[6650] = 1'b1;
assign COL[6651] = 1'b1;
assign COL[6652] = 1'b1;
assign COL[6653] = 1'b1;
assign COL[6654] = 1'b1;
assign COL[6655] = 1'b0;
assign COL[6656] = 1'b0;
assign COL[6657] = 1'b0;
assign COL[6658] = 1'b0;
assign COL[6659] = 1'b0;
assign COL[6660] = 1'b0;
assign COL[6661] = 1'b0;
assign COL[6662] = 1'b0;
assign COL[6663] = 1'b0;
assign COL[6664] = 1'b0;
assign COL[6665] = 1'b0;
assign COL[6666] = 1'b0;
assign COL[6667] = 1'b0;
assign COL[6668] = 1'b0;
assign COL[6669] = 1'b0;
assign COL[6670] = 1'b0;
assign COL[6671] = 1'b0;
assign COL[6672] = 1'b0;
assign COL[6673] = 1'b0;
assign COL[6674] = 1'b0;
assign COL[6675] = 1'b0;
assign COL[6676] = 1'b0;
assign COL[6677] = 1'b0;
assign COL[6678] = 1'b0;
assign COL[6679] = 1'b0;
assign COL[6680] = 1'b0;
assign COL[6681] = 1'b0;
assign COL[6682] = 1'b0;
assign COL[6683] = 1'b0;
assign COL[6684] = 1'b0;
assign COL[6685] = 1'b0;
assign COL[6686] = 1'b0;
assign COL[6687] = 1'b0;
assign COL[6688] = 1'b0;
assign COL[6689] = 1'b0;
assign COL[6690] = 1'b0;
assign COL[6691] = 1'b0;
assign COL[6692] = 1'b0;
assign COL[6693] = 1'b0;
assign COL[6694] = 1'b0;
assign COL[6695] = 1'b0;
assign COL[6696] = 1'b0;
assign COL[6697] = 1'b0;
assign COL[6698] = 1'b0;
assign COL[6699] = 1'b0;
assign COL[6700] = 1'b0;
assign COL[6701] = 1'b0;
assign COL[6702] = 1'b0;
assign COL[6703] = 1'b0;
assign COL[6704] = 1'b0;
assign COL[6705] = 1'b0;
assign COL[6706] = 1'b0;
assign COL[6707] = 1'b0;
assign COL[6708] = 1'b0;
assign COL[6709] = 1'b0;
assign COL[6710] = 1'b0;
assign COL[6711] = 1'b0;
assign COL[6712] = 1'b0;
assign COL[6713] = 1'b0;
assign COL[6714] = 1'b0;
assign COL[6715] = 1'b0;
assign COL[6716] = 1'b0;
assign COL[6717] = 1'b0;
assign COL[6718] = 1'b0;
assign COL[6719] = 1'b0;
assign COL[6720] = 1'b0;
assign COL[6721] = 1'b1;
assign COL[6722] = 1'b1;
assign COL[6723] = 1'b1;
assign COL[6724] = 1'b1;
assign COL[6725] = 1'b1;
assign COL[6726] = 1'b0;
assign COL[6727] = 1'b0;
assign COL[6728] = 1'b0;
assign COL[6729] = 1'b0;
assign COL[6730] = 1'b0;
assign COL[6731] = 1'b0;
assign COL[6732] = 1'b0;
assign COL[6733] = 1'b0;
assign COL[6734] = 1'b0;
assign COL[6735] = 1'b0;
assign COL[6736] = 1'b1;
assign COL[6737] = 1'b1;
assign COL[6738] = 1'b1;
assign COL[6739] = 1'b1;
assign COL[6740] = 1'b0;
assign COL[6741] = 1'b0;
assign COL[6742] = 1'b0;
assign COL[6743] = 1'b0;
assign COL[6744] = 1'b0;
assign COL[6745] = 1'b0;
assign COL[6746] = 1'b0;
assign COL[6747] = 1'b0;
assign COL[6748] = 1'b0;
assign COL[6749] = 1'b0;
assign COL[6750] = 1'b0;
assign COL[6751] = 1'b0;
assign COL[6752] = 1'b0;
assign COL[6753] = 1'b0;
assign COL[6754] = 1'b0;
assign COL[6755] = 1'b0;
assign COL[6756] = 1'b0;
assign COL[6757] = 1'b0;
assign COL[6758] = 1'b0;
assign COL[6759] = 1'b0;
assign COL[6760] = 1'b1;
assign COL[6761] = 1'b1;
assign COL[6762] = 1'b1;
assign COL[6763] = 1'b1;
assign COL[6764] = 1'b0;
assign COL[6765] = 1'b0;
assign COL[6766] = 1'b0;
assign COL[6767] = 1'b0;
assign COL[6768] = 1'b0;
assign COL[6769] = 1'b0;
assign COL[6770] = 1'b0;
assign COL[6771] = 1'b0;
assign COL[6772] = 1'b0;
assign COL[6773] = 1'b0;
assign COL[6774] = 1'b0;
assign COL[6775] = 1'b0;
assign COL[6776] = 1'b0;
assign COL[6777] = 1'b0;
assign COL[6778] = 1'b0;
assign COL[6779] = 1'b0;
assign COL[6780] = 1'b0;
assign COL[6781] = 1'b0;
assign COL[6782] = 1'b0;
assign COL[6783] = 1'b0;
assign COL[6784] = 1'b0;
assign COL[6785] = 1'b0;
assign COL[6786] = 1'b0;
assign COL[6787] = 1'b0;
assign COL[6788] = 1'b0;
assign COL[6789] = 1'b0;
assign COL[6790] = 1'b0;
assign COL[6791] = 1'b0;
assign COL[6792] = 1'b0;
assign COL[6793] = 1'b0;
assign COL[6794] = 1'b0;
assign COL[6795] = 1'b0;
assign COL[6796] = 1'b0;
assign COL[6797] = 1'b0;
assign COL[6798] = 1'b0;
assign COL[6799] = 1'b0;
assign COL[6800] = 1'b0;
assign COL[6801] = 1'b0;
assign COL[6802] = 1'b0;
assign COL[6803] = 1'b0;
assign COL[6804] = 1'b0;
assign COL[6805] = 1'b0;
assign COL[6806] = 1'b0;
assign COL[6807] = 1'b0;
assign COL[6808] = 1'b0;
assign COL[6809] = 1'b0;
assign COL[6810] = 1'b1;
assign COL[6811] = 1'b1;
assign COL[6812] = 1'b1;
assign COL[6813] = 1'b1;
assign COL[6814] = 1'b1;
assign COL[6815] = 1'b0;
assign COL[6816] = 1'b0;
assign COL[6817] = 1'b0;
assign COL[6818] = 1'b0;
assign COL[6819] = 1'b0;
assign COL[6820] = 1'b0;
assign COL[6821] = 1'b0;
assign COL[6822] = 1'b0;
assign COL[6823] = 1'b0;
assign COL[6824] = 1'b0;
assign COL[6825] = 1'b0;
assign COL[6826] = 1'b0;
assign COL[6827] = 1'b0;
assign COL[6828] = 1'b0;
assign COL[6829] = 1'b0;
assign COL[6830] = 1'b0;
assign COL[6831] = 1'b0;
assign COL[6832] = 1'b0;
assign COL[6833] = 1'b0;
assign COL[6834] = 1'b0;
assign COL[6835] = 1'b0;
assign COL[6836] = 1'b0;
assign COL[6837] = 1'b0;
assign COL[6838] = 1'b0;
assign COL[6839] = 1'b0;
assign COL[6840] = 1'b0;
assign COL[6841] = 1'b0;
assign COL[6842] = 1'b0;
assign COL[6843] = 1'b0;
assign COL[6844] = 1'b0;
assign COL[6845] = 1'b0;
assign COL[6846] = 1'b0;
assign COL[6847] = 1'b0;
assign COL[6848] = 1'b0;
assign COL[6849] = 1'b0;
assign COL[6850] = 1'b0;
assign COL[6851] = 1'b0;
assign COL[6852] = 1'b0;
assign COL[6853] = 1'b0;
assign COL[6854] = 1'b0;
assign COL[6855] = 1'b0;
assign COL[6856] = 1'b0;
assign COL[6857] = 1'b0;
assign COL[6858] = 1'b0;
assign COL[6859] = 1'b0;
assign COL[6860] = 1'b0;
assign COL[6861] = 1'b0;
assign COL[6862] = 1'b0;
assign COL[6863] = 1'b0;
assign COL[6864] = 1'b0;
assign COL[6865] = 1'b0;
assign COL[6866] = 1'b0;
assign COL[6867] = 1'b0;
assign COL[6868] = 1'b0;
assign COL[6869] = 1'b0;
assign COL[6870] = 1'b0;
assign COL[6871] = 1'b0;
assign COL[6872] = 1'b0;
assign COL[6873] = 1'b0;
assign COL[6874] = 1'b0;
assign COL[6875] = 1'b0;
assign COL[6876] = 1'b0;
assign COL[6877] = 1'b0;
assign COL[6878] = 1'b0;
assign COL[6879] = 1'b0;
assign COL[6880] = 1'b0;
assign COL[6881] = 1'b1;
assign COL[6882] = 1'b1;
assign COL[6883] = 1'b1;
assign COL[6884] = 1'b1;
assign COL[6885] = 1'b1;
assign COL[6886] = 1'b0;
assign COL[6887] = 1'b0;
assign COL[6888] = 1'b0;
assign COL[6889] = 1'b0;
assign COL[6890] = 1'b0;
assign COL[6891] = 1'b0;
assign COL[6892] = 1'b0;
assign COL[6893] = 1'b0;
assign COL[6894] = 1'b0;
assign COL[6895] = 1'b0;
assign COL[6896] = 1'b1;
assign COL[6897] = 1'b1;
assign COL[6898] = 1'b1;
assign COL[6899] = 1'b1;
assign COL[6900] = 1'b0;
assign COL[6901] = 1'b0;
assign COL[6902] = 1'b0;
assign COL[6903] = 1'b0;
assign COL[6904] = 1'b0;
assign COL[6905] = 1'b0;
assign COL[6906] = 1'b0;
assign COL[6907] = 1'b0;
assign COL[6908] = 1'b0;
assign COL[6909] = 1'b0;
assign COL[6910] = 1'b0;
assign COL[6911] = 1'b0;
assign COL[6912] = 1'b0;
assign COL[6913] = 1'b0;
assign COL[6914] = 1'b0;
assign COL[6915] = 1'b0;
assign COL[6916] = 1'b0;
assign COL[6917] = 1'b0;
assign COL[6918] = 1'b0;
assign COL[6919] = 1'b0;
assign COL[6920] = 1'b1;
assign COL[6921] = 1'b1;
assign COL[6922] = 1'b1;
assign COL[6923] = 1'b1;
assign COL[6924] = 1'b0;
assign COL[6925] = 1'b0;
assign COL[6926] = 1'b0;
assign COL[6927] = 1'b0;
assign COL[6928] = 1'b0;
assign COL[6929] = 1'b0;
assign COL[6930] = 1'b0;
assign COL[6931] = 1'b0;
assign COL[6932] = 1'b0;
assign COL[6933] = 1'b0;
assign COL[6934] = 1'b0;
assign COL[6935] = 1'b0;
assign COL[6936] = 1'b0;
assign COL[6937] = 1'b0;
assign COL[6938] = 1'b0;
assign COL[6939] = 1'b0;
assign COL[6940] = 1'b0;
assign COL[6941] = 1'b0;
assign COL[6942] = 1'b0;
assign COL[6943] = 1'b0;
assign COL[6944] = 1'b0;
assign COL[6945] = 1'b0;
assign COL[6946] = 1'b0;
assign COL[6947] = 1'b0;
assign COL[6948] = 1'b0;
assign COL[6949] = 1'b0;
assign COL[6950] = 1'b0;
assign COL[6951] = 1'b0;
assign COL[6952] = 1'b0;
assign COL[6953] = 1'b0;
assign COL[6954] = 1'b0;
assign COL[6955] = 1'b0;
assign COL[6956] = 1'b0;
assign COL[6957] = 1'b0;
assign COL[6958] = 1'b0;
assign COL[6959] = 1'b0;
assign COL[6960] = 1'b0;
assign COL[6961] = 1'b0;
assign COL[6962] = 1'b0;
assign COL[6963] = 1'b0;
assign COL[6964] = 1'b0;
assign COL[6965] = 1'b0;
assign COL[6966] = 1'b0;
assign COL[6967] = 1'b0;
assign COL[6968] = 1'b0;
assign COL[6969] = 1'b0;
assign COL[6970] = 1'b1;
assign COL[6971] = 1'b1;
assign COL[6972] = 1'b1;
assign COL[6973] = 1'b1;
assign COL[6974] = 1'b1;
assign COL[6975] = 1'b0;
assign COL[6976] = 1'b0;
assign COL[6977] = 1'b0;
assign COL[6978] = 1'b0;
assign COL[6979] = 1'b0;
assign COL[6980] = 1'b0;
assign COL[6981] = 1'b0;
assign COL[6982] = 1'b0;
assign COL[6983] = 1'b0;
assign COL[6984] = 1'b0;
assign COL[6985] = 1'b0;
assign COL[6986] = 1'b0;
assign COL[6987] = 1'b0;
assign COL[6988] = 1'b0;
assign COL[6989] = 1'b0;
assign COL[6990] = 1'b0;
assign COL[6991] = 1'b0;
assign COL[6992] = 1'b0;
assign COL[6993] = 1'b0;
assign COL[6994] = 1'b0;
assign COL[6995] = 1'b0;
assign COL[6996] = 1'b0;
assign COL[6997] = 1'b0;
assign COL[6998] = 1'b0;
assign COL[6999] = 1'b0;
assign COL[7000] = 1'b0;
assign COL[7001] = 1'b0;
assign COL[7002] = 1'b0;
assign COL[7003] = 1'b0;
assign COL[7004] = 1'b0;
assign COL[7005] = 1'b0;
assign COL[7006] = 1'b0;
assign COL[7007] = 1'b0;
assign COL[7008] = 1'b0;
assign COL[7009] = 1'b0;
assign COL[7010] = 1'b0;
assign COL[7011] = 1'b0;
assign COL[7012] = 1'b0;
assign COL[7013] = 1'b0;
assign COL[7014] = 1'b0;
assign COL[7015] = 1'b0;
assign COL[7016] = 1'b0;
assign COL[7017] = 1'b0;
assign COL[7018] = 1'b0;
assign COL[7019] = 1'b0;
assign COL[7020] = 1'b0;
assign COL[7021] = 1'b0;
assign COL[7022] = 1'b0;
assign COL[7023] = 1'b0;
assign COL[7024] = 1'b0;
assign COL[7025] = 1'b0;
assign COL[7026] = 1'b0;
assign COL[7027] = 1'b0;
assign COL[7028] = 1'b0;
assign COL[7029] = 1'b0;
assign COL[7030] = 1'b0;
assign COL[7031] = 1'b0;
assign COL[7032] = 1'b0;
assign COL[7033] = 1'b0;
assign COL[7034] = 1'b0;
assign COL[7035] = 1'b0;
assign COL[7036] = 1'b0;
assign COL[7037] = 1'b0;
assign COL[7038] = 1'b0;
assign COL[7039] = 1'b0;
assign COL[7040] = 1'b0;
assign COL[7041] = 1'b1;
assign COL[7042] = 1'b1;
assign COL[7043] = 1'b1;
assign COL[7044] = 1'b1;
assign COL[7045] = 1'b1;
assign COL[7046] = 1'b0;
assign COL[7047] = 1'b0;
assign COL[7048] = 1'b0;
assign COL[7049] = 1'b0;
assign COL[7050] = 1'b0;
assign COL[7051] = 1'b0;
assign COL[7052] = 1'b0;
assign COL[7053] = 1'b0;
assign COL[7054] = 1'b0;
assign COL[7055] = 1'b0;
assign COL[7056] = 1'b1;
assign COL[7057] = 1'b1;
assign COL[7058] = 1'b1;
assign COL[7059] = 1'b1;
assign COL[7060] = 1'b0;
assign COL[7061] = 1'b0;
assign COL[7062] = 1'b0;
assign COL[7063] = 1'b0;
assign COL[7064] = 1'b0;
assign COL[7065] = 1'b0;
assign COL[7066] = 1'b0;
assign COL[7067] = 1'b0;
assign COL[7068] = 1'b0;
assign COL[7069] = 1'b0;
assign COL[7070] = 1'b0;
assign COL[7071] = 1'b0;
assign COL[7072] = 1'b0;
assign COL[7073] = 1'b0;
assign COL[7074] = 1'b0;
assign COL[7075] = 1'b0;
assign COL[7076] = 1'b0;
assign COL[7077] = 1'b0;
assign COL[7078] = 1'b0;
assign COL[7079] = 1'b0;
assign COL[7080] = 1'b1;
assign COL[7081] = 1'b1;
assign COL[7082] = 1'b1;
assign COL[7083] = 1'b1;
assign COL[7084] = 1'b0;
assign COL[7085] = 1'b0;
assign COL[7086] = 1'b0;
assign COL[7087] = 1'b0;
assign COL[7088] = 1'b0;
assign COL[7089] = 1'b0;
assign COL[7090] = 1'b0;
assign COL[7091] = 1'b0;
assign COL[7092] = 1'b0;
assign COL[7093] = 1'b0;
assign COL[7094] = 1'b0;
assign COL[7095] = 1'b0;
assign COL[7096] = 1'b0;
assign COL[7097] = 1'b0;
assign COL[7098] = 1'b0;
assign COL[7099] = 1'b0;
assign COL[7100] = 1'b0;
assign COL[7101] = 1'b0;
assign COL[7102] = 1'b0;
assign COL[7103] = 1'b0;
assign COL[7104] = 1'b0;
assign COL[7105] = 1'b0;
assign COL[7106] = 1'b0;
assign COL[7107] = 1'b0;
assign COL[7108] = 1'b0;
assign COL[7109] = 1'b0;
assign COL[7110] = 1'b0;
assign COL[7111] = 1'b0;
assign COL[7112] = 1'b0;
assign COL[7113] = 1'b0;
assign COL[7114] = 1'b0;
assign COL[7115] = 1'b0;
assign COL[7116] = 1'b0;
assign COL[7117] = 1'b0;
assign COL[7118] = 1'b0;
assign COL[7119] = 1'b0;
assign COL[7120] = 1'b0;
assign COL[7121] = 1'b0;
assign COL[7122] = 1'b0;
assign COL[7123] = 1'b0;
assign COL[7124] = 1'b0;
assign COL[7125] = 1'b0;
assign COL[7126] = 1'b0;
assign COL[7127] = 1'b0;
assign COL[7128] = 1'b0;
assign COL[7129] = 1'b0;
assign COL[7130] = 1'b1;
assign COL[7131] = 1'b1;
assign COL[7132] = 1'b1;
assign COL[7133] = 1'b1;
assign COL[7134] = 1'b1;
assign COL[7135] = 1'b0;
assign COL[7136] = 1'b0;
assign COL[7137] = 1'b0;
assign COL[7138] = 1'b0;
assign COL[7139] = 1'b0;
assign COL[7140] = 1'b0;
assign COL[7141] = 1'b0;
assign COL[7142] = 1'b0;
assign COL[7143] = 1'b0;
assign COL[7144] = 1'b0;
assign COL[7145] = 1'b0;
assign COL[7146] = 1'b0;
assign COL[7147] = 1'b0;
assign COL[7148] = 1'b0;
assign COL[7149] = 1'b0;
assign COL[7150] = 1'b0;
assign COL[7151] = 1'b0;
assign COL[7152] = 1'b0;
assign COL[7153] = 1'b0;
assign COL[7154] = 1'b0;
assign COL[7155] = 1'b0;
assign COL[7156] = 1'b0;
assign COL[7157] = 1'b0;
assign COL[7158] = 1'b0;
assign COL[7159] = 1'b0;
assign COL[7160] = 1'b0;
assign COL[7161] = 1'b0;
assign COL[7162] = 1'b0;
assign COL[7163] = 1'b0;
assign COL[7164] = 1'b0;
assign COL[7165] = 1'b0;
assign COL[7166] = 1'b0;
assign COL[7167] = 1'b0;
assign COL[7168] = 1'b0;
assign COL[7169] = 1'b0;
assign COL[7170] = 1'b0;
assign COL[7171] = 1'b0;
assign COL[7172] = 1'b0;
assign COL[7173] = 1'b0;
assign COL[7174] = 1'b0;
assign COL[7175] = 1'b0;
assign COL[7176] = 1'b0;
assign COL[7177] = 1'b0;
assign COL[7178] = 1'b0;
assign COL[7179] = 1'b0;
assign COL[7180] = 1'b0;
assign COL[7181] = 1'b0;
assign COL[7182] = 1'b0;
assign COL[7183] = 1'b0;
assign COL[7184] = 1'b0;
assign COL[7185] = 1'b0;
assign COL[7186] = 1'b0;
assign COL[7187] = 1'b0;
assign COL[7188] = 1'b0;
assign COL[7189] = 1'b0;
assign COL[7190] = 1'b0;
assign COL[7191] = 1'b0;
assign COL[7192] = 1'b0;
assign COL[7193] = 1'b0;
assign COL[7194] = 1'b0;
assign COL[7195] = 1'b0;
assign COL[7196] = 1'b0;
assign COL[7197] = 1'b0;
assign COL[7198] = 1'b0;
assign COL[7199] = 1'b0;
assign COL[7200] = 1'b0;
assign COL[7201] = 1'b1;
assign COL[7202] = 1'b1;
assign COL[7203] = 1'b1;
assign COL[7204] = 1'b1;
assign COL[7205] = 1'b1;
assign COL[7206] = 1'b0;
assign COL[7207] = 1'b0;
assign COL[7208] = 1'b0;
assign COL[7209] = 1'b0;
assign COL[7210] = 1'b0;
assign COL[7211] = 1'b0;
assign COL[7212] = 1'b0;
assign COL[7213] = 1'b0;
assign COL[7214] = 1'b0;
assign COL[7215] = 1'b0;
assign COL[7216] = 1'b1;
assign COL[7217] = 1'b1;
assign COL[7218] = 1'b1;
assign COL[7219] = 1'b1;
assign COL[7220] = 1'b0;
assign COL[7221] = 1'b0;
assign COL[7222] = 1'b0;
assign COL[7223] = 1'b0;
assign COL[7224] = 1'b0;
assign COL[7225] = 1'b0;
assign COL[7226] = 1'b0;
assign COL[7227] = 1'b0;
assign COL[7228] = 1'b0;
assign COL[7229] = 1'b0;
assign COL[7230] = 1'b0;
assign COL[7231] = 1'b0;
assign COL[7232] = 1'b0;
assign COL[7233] = 1'b0;
assign COL[7234] = 1'b0;
assign COL[7235] = 1'b0;
assign COL[7236] = 1'b0;
assign COL[7237] = 1'b0;
assign COL[7238] = 1'b0;
assign COL[7239] = 1'b0;
assign COL[7240] = 1'b1;
assign COL[7241] = 1'b1;
assign COL[7242] = 1'b1;
assign COL[7243] = 1'b1;
assign COL[7244] = 1'b0;
assign COL[7245] = 1'b0;
assign COL[7246] = 1'b0;
assign COL[7247] = 1'b0;
assign COL[7248] = 1'b0;
assign COL[7249] = 1'b0;
assign COL[7250] = 1'b0;
assign COL[7251] = 1'b0;
assign COL[7252] = 1'b0;
assign COL[7253] = 1'b0;
assign COL[7254] = 1'b0;
assign COL[7255] = 1'b0;
assign COL[7256] = 1'b0;
assign COL[7257] = 1'b0;
assign COL[7258] = 1'b0;
assign COL[7259] = 1'b0;
assign COL[7260] = 1'b0;
assign COL[7261] = 1'b0;
assign COL[7262] = 1'b0;
assign COL[7263] = 1'b0;
assign COL[7264] = 1'b0;
assign COL[7265] = 1'b0;
assign COL[7266] = 1'b0;
assign COL[7267] = 1'b0;
assign COL[7268] = 1'b0;
assign COL[7269] = 1'b0;
assign COL[7270] = 1'b0;
assign COL[7271] = 1'b0;
assign COL[7272] = 1'b0;
assign COL[7273] = 1'b0;
assign COL[7274] = 1'b0;
assign COL[7275] = 1'b0;
assign COL[7276] = 1'b0;
assign COL[7277] = 1'b0;
assign COL[7278] = 1'b0;
assign COL[7279] = 1'b0;
assign COL[7280] = 1'b0;
assign COL[7281] = 1'b0;
assign COL[7282] = 1'b0;
assign COL[7283] = 1'b0;
assign COL[7284] = 1'b0;
assign COL[7285] = 1'b0;
assign COL[7286] = 1'b0;
assign COL[7287] = 1'b0;
assign COL[7288] = 1'b0;
assign COL[7289] = 1'b0;
assign COL[7290] = 1'b1;
assign COL[7291] = 1'b1;
assign COL[7292] = 1'b1;
assign COL[7293] = 1'b1;
assign COL[7294] = 1'b1;
assign COL[7295] = 1'b0;
assign COL[7296] = 1'b0;
assign COL[7297] = 1'b0;
assign COL[7298] = 1'b0;
assign COL[7299] = 1'b0;
assign COL[7300] = 1'b0;
assign COL[7301] = 1'b0;
assign COL[7302] = 1'b0;
assign COL[7303] = 1'b0;
assign COL[7304] = 1'b0;
assign COL[7305] = 1'b0;
assign COL[7306] = 1'b0;
assign COL[7307] = 1'b0;
assign COL[7308] = 1'b0;
assign COL[7309] = 1'b0;
assign COL[7310] = 1'b0;
assign COL[7311] = 1'b0;
assign COL[7312] = 1'b0;
assign COL[7313] = 1'b0;
assign COL[7314] = 1'b0;
assign COL[7315] = 1'b0;
assign COL[7316] = 1'b0;
assign COL[7317] = 1'b0;
assign COL[7318] = 1'b0;
assign COL[7319] = 1'b0;
assign COL[7320] = 1'b0;
assign COL[7321] = 1'b0;
assign COL[7322] = 1'b0;
assign COL[7323] = 1'b0;
assign COL[7324] = 1'b0;
assign COL[7325] = 1'b0;
assign COL[7326] = 1'b0;
assign COL[7327] = 1'b0;
assign COL[7328] = 1'b0;
assign COL[7329] = 1'b0;
assign COL[7330] = 1'b0;
assign COL[7331] = 1'b0;
assign COL[7332] = 1'b0;
assign COL[7333] = 1'b0;
assign COL[7334] = 1'b0;
assign COL[7335] = 1'b0;
assign COL[7336] = 1'b0;
assign COL[7337] = 1'b0;
assign COL[7338] = 1'b0;
assign COL[7339] = 1'b0;
assign COL[7340] = 1'b0;
assign COL[7341] = 1'b0;
assign COL[7342] = 1'b0;
assign COL[7343] = 1'b0;
assign COL[7344] = 1'b0;
assign COL[7345] = 1'b0;
assign COL[7346] = 1'b0;
assign COL[7347] = 1'b0;
assign COL[7348] = 1'b0;
assign COL[7349] = 1'b0;
assign COL[7350] = 1'b0;
assign COL[7351] = 1'b0;
assign COL[7352] = 1'b0;
assign COL[7353] = 1'b0;
assign COL[7354] = 1'b0;
assign COL[7355] = 1'b0;
assign COL[7356] = 1'b0;
assign COL[7357] = 1'b0;
assign COL[7358] = 1'b0;
assign COL[7359] = 1'b0;
assign COL[7360] = 1'b0;
assign COL[7361] = 1'b1;
assign COL[7362] = 1'b1;
assign COL[7363] = 1'b1;
assign COL[7364] = 1'b1;
assign COL[7365] = 1'b1;
assign COL[7366] = 1'b0;
assign COL[7367] = 1'b0;
assign COL[7368] = 1'b0;
assign COL[7369] = 1'b0;
assign COL[7370] = 1'b0;
assign COL[7371] = 1'b0;
assign COL[7372] = 1'b0;
assign COL[7373] = 1'b0;
assign COL[7374] = 1'b0;
assign COL[7375] = 1'b0;
assign COL[7376] = 1'b1;
assign COL[7377] = 1'b1;
assign COL[7378] = 1'b1;
assign COL[7379] = 1'b1;
assign COL[7380] = 1'b0;
assign COL[7381] = 1'b0;
assign COL[7382] = 1'b0;
assign COL[7383] = 1'b0;
assign COL[7384] = 1'b0;
assign COL[7385] = 1'b0;
assign COL[7386] = 1'b0;
assign COL[7387] = 1'b0;
assign COL[7388] = 1'b0;
assign COL[7389] = 1'b0;
assign COL[7390] = 1'b0;
assign COL[7391] = 1'b0;
assign COL[7392] = 1'b0;
assign COL[7393] = 1'b0;
assign COL[7394] = 1'b0;
assign COL[7395] = 1'b0;
assign COL[7396] = 1'b0;
assign COL[7397] = 1'b0;
assign COL[7398] = 1'b0;
assign COL[7399] = 1'b0;
assign COL[7400] = 1'b1;
assign COL[7401] = 1'b1;
assign COL[7402] = 1'b1;
assign COL[7403] = 1'b1;
assign COL[7404] = 1'b0;
assign COL[7405] = 1'b0;
assign COL[7406] = 1'b0;
assign COL[7407] = 1'b0;
assign COL[7408] = 1'b0;
assign COL[7409] = 1'b0;
assign COL[7410] = 1'b0;
assign COL[7411] = 1'b0;
assign COL[7412] = 1'b0;
assign COL[7413] = 1'b0;
assign COL[7414] = 1'b0;
assign COL[7415] = 1'b0;
assign COL[7416] = 1'b0;
assign COL[7417] = 1'b0;
assign COL[7418] = 1'b0;
assign COL[7419] = 1'b0;
assign COL[7420] = 1'b0;
assign COL[7421] = 1'b0;
assign COL[7422] = 1'b0;
assign COL[7423] = 1'b0;
assign COL[7424] = 1'b0;
assign COL[7425] = 1'b0;
assign COL[7426] = 1'b0;
assign COL[7427] = 1'b0;
assign COL[7428] = 1'b0;
assign COL[7429] = 1'b0;
assign COL[7430] = 1'b0;
assign COL[7431] = 1'b0;
assign COL[7432] = 1'b0;
assign COL[7433] = 1'b0;
assign COL[7434] = 1'b0;
assign COL[7435] = 1'b0;
assign COL[7436] = 1'b0;
assign COL[7437] = 1'b0;
assign COL[7438] = 1'b0;
assign COL[7439] = 1'b0;
assign COL[7440] = 1'b0;
assign COL[7441] = 1'b0;
assign COL[7442] = 1'b0;
assign COL[7443] = 1'b0;
assign COL[7444] = 1'b0;
assign COL[7445] = 1'b0;
assign COL[7446] = 1'b0;
assign COL[7447] = 1'b0;
assign COL[7448] = 1'b0;
assign COL[7449] = 1'b0;
assign COL[7450] = 1'b1;
assign COL[7451] = 1'b1;
assign COL[7452] = 1'b1;
assign COL[7453] = 1'b1;
assign COL[7454] = 1'b1;
assign COL[7455] = 1'b0;
assign COL[7456] = 1'b0;
assign COL[7457] = 1'b0;
assign COL[7458] = 1'b0;
assign COL[7459] = 1'b0;
assign COL[7460] = 1'b0;
assign COL[7461] = 1'b0;
assign COL[7462] = 1'b0;
assign COL[7463] = 1'b0;
assign COL[7464] = 1'b0;
assign COL[7465] = 1'b0;
assign COL[7466] = 1'b0;
assign COL[7467] = 1'b0;
assign COL[7468] = 1'b0;
assign COL[7469] = 1'b0;
assign COL[7470] = 1'b0;
assign COL[7471] = 1'b0;
assign COL[7472] = 1'b0;
assign COL[7473] = 1'b0;
assign COL[7474] = 1'b0;
assign COL[7475] = 1'b0;
assign COL[7476] = 1'b0;
assign COL[7477] = 1'b0;
assign COL[7478] = 1'b0;
assign COL[7479] = 1'b0;
assign COL[7480] = 1'b0;
assign COL[7481] = 1'b0;
assign COL[7482] = 1'b0;
assign COL[7483] = 1'b0;
assign COL[7484] = 1'b0;
assign COL[7485] = 1'b0;
assign COL[7486] = 1'b0;
assign COL[7487] = 1'b0;
assign COL[7488] = 1'b0;
assign COL[7489] = 1'b0;
assign COL[7490] = 1'b0;
assign COL[7491] = 1'b0;
assign COL[7492] = 1'b0;
assign COL[7493] = 1'b0;
assign COL[7494] = 1'b0;
assign COL[7495] = 1'b0;
assign COL[7496] = 1'b0;
assign COL[7497] = 1'b0;
assign COL[7498] = 1'b0;
assign COL[7499] = 1'b0;
assign COL[7500] = 1'b0;
assign COL[7501] = 1'b0;
assign COL[7502] = 1'b0;
assign COL[7503] = 1'b0;
assign COL[7504] = 1'b0;
assign COL[7505] = 1'b0;
assign COL[7506] = 1'b0;
assign COL[7507] = 1'b0;
assign COL[7508] = 1'b0;
assign COL[7509] = 1'b0;
assign COL[7510] = 1'b0;
assign COL[7511] = 1'b0;
assign COL[7512] = 1'b0;
assign COL[7513] = 1'b0;
assign COL[7514] = 1'b0;
assign COL[7515] = 1'b0;
assign COL[7516] = 1'b0;
assign COL[7517] = 1'b0;
assign COL[7518] = 1'b0;
assign COL[7519] = 1'b0;
assign COL[7520] = 1'b0;
assign COL[7521] = 1'b1;
assign COL[7522] = 1'b1;
assign COL[7523] = 1'b1;
assign COL[7524] = 1'b1;
assign COL[7525] = 1'b1;
assign COL[7526] = 1'b0;
assign COL[7527] = 1'b0;
assign COL[7528] = 1'b0;
assign COL[7529] = 1'b0;
assign COL[7530] = 1'b0;
assign COL[7531] = 1'b0;
assign COL[7532] = 1'b0;
assign COL[7533] = 1'b0;
assign COL[7534] = 1'b0;
assign COL[7535] = 1'b0;
assign COL[7536] = 1'b1;
assign COL[7537] = 1'b1;
assign COL[7538] = 1'b1;
assign COL[7539] = 1'b1;
assign COL[7540] = 1'b1;
assign COL[7541] = 1'b1;
assign COL[7542] = 1'b1;
assign COL[7543] = 1'b1;
assign COL[7544] = 1'b1;
assign COL[7545] = 1'b1;
assign COL[7546] = 1'b1;
assign COL[7547] = 1'b1;
assign COL[7548] = 1'b1;
assign COL[7549] = 1'b1;
assign COL[7550] = 1'b1;
assign COL[7551] = 1'b1;
assign COL[7552] = 1'b1;
assign COL[7553] = 1'b1;
assign COL[7554] = 1'b1;
assign COL[7555] = 1'b1;
assign COL[7556] = 1'b1;
assign COL[7557] = 1'b1;
assign COL[7558] = 1'b1;
assign COL[7559] = 1'b1;
assign COL[7560] = 1'b1;
assign COL[7561] = 1'b1;
assign COL[7562] = 1'b1;
assign COL[7563] = 1'b1;
assign COL[7564] = 1'b1;
assign COL[7565] = 1'b1;
assign COL[7566] = 1'b1;
assign COL[7567] = 1'b1;
assign COL[7568] = 1'b1;
assign COL[7569] = 1'b1;
assign COL[7570] = 1'b1;
assign COL[7571] = 1'b1;
assign COL[7572] = 1'b1;
assign COL[7573] = 1'b1;
assign COL[7574] = 1'b1;
assign COL[7575] = 1'b1;
assign COL[7576] = 1'b1;
assign COL[7577] = 1'b1;
assign COL[7578] = 1'b1;
assign COL[7579] = 1'b1;
assign COL[7580] = 1'b1;
assign COL[7581] = 1'b1;
assign COL[7582] = 1'b0;
assign COL[7583] = 1'b0;
assign COL[7584] = 1'b0;
assign COL[7585] = 1'b0;
assign COL[7586] = 1'b0;
assign COL[7587] = 1'b0;
assign COL[7588] = 1'b0;
assign COL[7589] = 1'b0;
assign COL[7590] = 1'b0;
assign COL[7591] = 1'b0;
assign COL[7592] = 1'b0;
assign COL[7593] = 1'b0;
assign COL[7594] = 1'b0;
assign COL[7595] = 1'b0;
assign COL[7596] = 1'b0;
assign COL[7597] = 1'b0;
assign COL[7598] = 1'b0;
assign COL[7599] = 1'b0;
assign COL[7600] = 1'b0;
assign COL[7601] = 1'b0;
assign COL[7602] = 1'b0;
assign COL[7603] = 1'b0;
assign COL[7604] = 1'b0;
assign COL[7605] = 1'b0;
assign COL[7606] = 1'b0;
assign COL[7607] = 1'b0;
assign COL[7608] = 1'b0;
assign COL[7609] = 1'b0;
assign COL[7610] = 1'b1;
assign COL[7611] = 1'b1;
assign COL[7612] = 1'b1;
assign COL[7613] = 1'b1;
assign COL[7614] = 1'b1;
assign COL[7615] = 1'b0;
assign COL[7616] = 1'b0;
assign COL[7617] = 1'b0;
assign COL[7618] = 1'b0;
assign COL[7619] = 1'b0;
assign COL[7620] = 1'b0;
assign COL[7621] = 1'b0;
assign COL[7622] = 1'b0;
assign COL[7623] = 1'b0;
assign COL[7624] = 1'b0;
assign COL[7625] = 1'b0;
assign COL[7626] = 1'b0;
assign COL[7627] = 1'b0;
assign COL[7628] = 1'b0;
assign COL[7629] = 1'b0;
assign COL[7630] = 1'b0;
assign COL[7631] = 1'b0;
assign COL[7632] = 1'b0;
assign COL[7633] = 1'b0;
assign COL[7634] = 1'b0;
assign COL[7635] = 1'b0;
assign COL[7636] = 1'b0;
assign COL[7637] = 1'b0;
assign COL[7638] = 1'b0;
assign COL[7639] = 1'b0;
assign COL[7640] = 1'b0;
assign COL[7641] = 1'b0;
assign COL[7642] = 1'b0;
assign COL[7643] = 1'b0;
assign COL[7644] = 1'b0;
assign COL[7645] = 1'b0;
assign COL[7646] = 1'b0;
assign COL[7647] = 1'b0;
assign COL[7648] = 1'b0;
assign COL[7649] = 1'b0;
assign COL[7650] = 1'b0;
assign COL[7651] = 1'b0;
assign COL[7652] = 1'b0;
assign COL[7653] = 1'b0;
assign COL[7654] = 1'b0;
assign COL[7655] = 1'b0;
assign COL[7656] = 1'b0;
assign COL[7657] = 1'b0;
assign COL[7658] = 1'b0;
assign COL[7659] = 1'b0;
assign COL[7660] = 1'b0;
assign COL[7661] = 1'b0;
assign COL[7662] = 1'b0;
assign COL[7663] = 1'b0;
assign COL[7664] = 1'b0;
assign COL[7665] = 1'b0;
assign COL[7666] = 1'b0;
assign COL[7667] = 1'b0;
assign COL[7668] = 1'b0;
assign COL[7669] = 1'b0;
assign COL[7670] = 1'b0;
assign COL[7671] = 1'b0;
assign COL[7672] = 1'b0;
assign COL[7673] = 1'b0;
assign COL[7674] = 1'b0;
assign COL[7675] = 1'b0;
assign COL[7676] = 1'b0;
assign COL[7677] = 1'b0;
assign COL[7678] = 1'b0;
assign COL[7679] = 1'b0;
assign COL[7680] = 1'b0;
assign COL[7681] = 1'b1;
assign COL[7682] = 1'b1;
assign COL[7683] = 1'b1;
assign COL[7684] = 1'b1;
assign COL[7685] = 1'b1;
assign COL[7686] = 1'b0;
assign COL[7687] = 1'b0;
assign COL[7688] = 1'b0;
assign COL[7689] = 1'b0;
assign COL[7690] = 1'b0;
assign COL[7691] = 1'b0;
assign COL[7692] = 1'b0;
assign COL[7693] = 1'b0;
assign COL[7694] = 1'b0;
assign COL[7695] = 1'b0;
assign COL[7696] = 1'b1;
assign COL[7697] = 1'b1;
assign COL[7698] = 1'b1;
assign COL[7699] = 1'b1;
assign COL[7700] = 1'b1;
assign COL[7701] = 1'b1;
assign COL[7702] = 1'b1;
assign COL[7703] = 1'b1;
assign COL[7704] = 1'b1;
assign COL[7705] = 1'b1;
assign COL[7706] = 1'b1;
assign COL[7707] = 1'b1;
assign COL[7708] = 1'b1;
assign COL[7709] = 1'b1;
assign COL[7710] = 1'b1;
assign COL[7711] = 1'b1;
assign COL[7712] = 1'b1;
assign COL[7713] = 1'b1;
assign COL[7714] = 1'b1;
assign COL[7715] = 1'b1;
assign COL[7716] = 1'b1;
assign COL[7717] = 1'b1;
assign COL[7718] = 1'b1;
assign COL[7719] = 1'b1;
assign COL[7720] = 1'b1;
assign COL[7721] = 1'b1;
assign COL[7722] = 1'b1;
assign COL[7723] = 1'b1;
assign COL[7724] = 1'b1;
assign COL[7725] = 1'b1;
assign COL[7726] = 1'b1;
assign COL[7727] = 1'b1;
assign COL[7728] = 1'b1;
assign COL[7729] = 1'b1;
assign COL[7730] = 1'b1;
assign COL[7731] = 1'b1;
assign COL[7732] = 1'b1;
assign COL[7733] = 1'b1;
assign COL[7734] = 1'b1;
assign COL[7735] = 1'b1;
assign COL[7736] = 1'b1;
assign COL[7737] = 1'b1;
assign COL[7738] = 1'b1;
assign COL[7739] = 1'b1;
assign COL[7740] = 1'b1;
assign COL[7741] = 1'b1;
assign COL[7742] = 1'b0;
assign COL[7743] = 1'b0;
assign COL[7744] = 1'b0;
assign COL[7745] = 1'b0;
assign COL[7746] = 1'b0;
assign COL[7747] = 1'b0;
assign COL[7748] = 1'b0;
assign COL[7749] = 1'b0;
assign COL[7750] = 1'b0;
assign COL[7751] = 1'b0;
assign COL[7752] = 1'b0;
assign COL[7753] = 1'b0;
assign COL[7754] = 1'b0;
assign COL[7755] = 1'b0;
assign COL[7756] = 1'b0;
assign COL[7757] = 1'b0;
assign COL[7758] = 1'b0;
assign COL[7759] = 1'b0;
assign COL[7760] = 1'b0;
assign COL[7761] = 1'b0;
assign COL[7762] = 1'b0;
assign COL[7763] = 1'b0;
assign COL[7764] = 1'b0;
assign COL[7765] = 1'b0;
assign COL[7766] = 1'b0;
assign COL[7767] = 1'b0;
assign COL[7768] = 1'b0;
assign COL[7769] = 1'b0;
assign COL[7770] = 1'b1;
assign COL[7771] = 1'b1;
assign COL[7772] = 1'b1;
assign COL[7773] = 1'b1;
assign COL[7774] = 1'b1;
assign COL[7775] = 1'b0;
assign COL[7776] = 1'b0;
assign COL[7777] = 1'b0;
assign COL[7778] = 1'b0;
assign COL[7779] = 1'b0;
assign COL[7780] = 1'b0;
assign COL[7781] = 1'b0;
assign COL[7782] = 1'b0;
assign COL[7783] = 1'b0;
assign COL[7784] = 1'b0;
assign COL[7785] = 1'b0;
assign COL[7786] = 1'b0;
assign COL[7787] = 1'b0;
assign COL[7788] = 1'b0;
assign COL[7789] = 1'b0;
assign COL[7790] = 1'b0;
assign COL[7791] = 1'b0;
assign COL[7792] = 1'b0;
assign COL[7793] = 1'b0;
assign COL[7794] = 1'b0;
assign COL[7795] = 1'b0;
assign COL[7796] = 1'b0;
assign COL[7797] = 1'b0;
assign COL[7798] = 1'b0;
assign COL[7799] = 1'b0;
assign COL[7800] = 1'b0;
assign COL[7801] = 1'b0;
assign COL[7802] = 1'b0;
assign COL[7803] = 1'b0;
assign COL[7804] = 1'b0;
assign COL[7805] = 1'b0;
assign COL[7806] = 1'b0;
assign COL[7807] = 1'b0;
assign COL[7808] = 1'b0;
assign COL[7809] = 1'b0;
assign COL[7810] = 1'b0;
assign COL[7811] = 1'b0;
assign COL[7812] = 1'b0;
assign COL[7813] = 1'b0;
assign COL[7814] = 1'b0;
assign COL[7815] = 1'b0;
assign COL[7816] = 1'b0;
assign COL[7817] = 1'b0;
assign COL[7818] = 1'b0;
assign COL[7819] = 1'b0;
assign COL[7820] = 1'b0;
assign COL[7821] = 1'b0;
assign COL[7822] = 1'b0;
assign COL[7823] = 1'b0;
assign COL[7824] = 1'b0;
assign COL[7825] = 1'b0;
assign COL[7826] = 1'b0;
assign COL[7827] = 1'b0;
assign COL[7828] = 1'b0;
assign COL[7829] = 1'b0;
assign COL[7830] = 1'b0;
assign COL[7831] = 1'b0;
assign COL[7832] = 1'b0;
assign COL[7833] = 1'b0;
assign COL[7834] = 1'b0;
assign COL[7835] = 1'b0;
assign COL[7836] = 1'b0;
assign COL[7837] = 1'b0;
assign COL[7838] = 1'b0;
assign COL[7839] = 1'b0;
assign COL[7840] = 1'b0;
assign COL[7841] = 1'b1;
assign COL[7842] = 1'b1;
assign COL[7843] = 1'b1;
assign COL[7844] = 1'b1;
assign COL[7845] = 1'b1;
assign COL[7846] = 1'b0;
assign COL[7847] = 1'b0;
assign COL[7848] = 1'b0;
assign COL[7849] = 1'b0;
assign COL[7850] = 1'b0;
assign COL[7851] = 1'b0;
assign COL[7852] = 1'b0;
assign COL[7853] = 1'b0;
assign COL[7854] = 1'b0;
assign COL[7855] = 1'b0;
assign COL[7856] = 1'b1;
assign COL[7857] = 1'b1;
assign COL[7858] = 1'b1;
assign COL[7859] = 1'b1;
assign COL[7860] = 1'b1;
assign COL[7861] = 1'b1;
assign COL[7862] = 1'b1;
assign COL[7863] = 1'b1;
assign COL[7864] = 1'b1;
assign COL[7865] = 1'b1;
assign COL[7866] = 1'b1;
assign COL[7867] = 1'b1;
assign COL[7868] = 1'b1;
assign COL[7869] = 1'b1;
assign COL[7870] = 1'b1;
assign COL[7871] = 1'b1;
assign COL[7872] = 1'b1;
assign COL[7873] = 1'b1;
assign COL[7874] = 1'b1;
assign COL[7875] = 1'b1;
assign COL[7876] = 1'b1;
assign COL[7877] = 1'b1;
assign COL[7878] = 1'b1;
assign COL[7879] = 1'b1;
assign COL[7880] = 1'b1;
assign COL[7881] = 1'b1;
assign COL[7882] = 1'b1;
assign COL[7883] = 1'b1;
assign COL[7884] = 1'b1;
assign COL[7885] = 1'b1;
assign COL[7886] = 1'b1;
assign COL[7887] = 1'b1;
assign COL[7888] = 1'b1;
assign COL[7889] = 1'b1;
assign COL[7890] = 1'b1;
assign COL[7891] = 1'b1;
assign COL[7892] = 1'b1;
assign COL[7893] = 1'b1;
assign COL[7894] = 1'b1;
assign COL[7895] = 1'b1;
assign COL[7896] = 1'b1;
assign COL[7897] = 1'b1;
assign COL[7898] = 1'b1;
assign COL[7899] = 1'b1;
assign COL[7900] = 1'b1;
assign COL[7901] = 1'b1;
assign COL[7902] = 1'b0;
assign COL[7903] = 1'b0;
assign COL[7904] = 1'b0;
assign COL[7905] = 1'b0;
assign COL[7906] = 1'b0;
assign COL[7907] = 1'b0;
assign COL[7908] = 1'b0;
assign COL[7909] = 1'b0;
assign COL[7910] = 1'b1;
assign COL[7911] = 1'b1;
assign COL[7912] = 1'b1;
assign COL[7913] = 1'b1;
assign COL[7914] = 1'b1;
assign COL[7915] = 1'b0;
assign COL[7916] = 1'b0;
assign COL[7917] = 1'b0;
assign COL[7918] = 1'b0;
assign COL[7919] = 1'b0;
assign COL[7920] = 1'b0;
assign COL[7921] = 1'b0;
assign COL[7922] = 1'b0;
assign COL[7923] = 1'b0;
assign COL[7924] = 1'b0;
assign COL[7925] = 1'b0;
assign COL[7926] = 1'b0;
assign COL[7927] = 1'b0;
assign COL[7928] = 1'b0;
assign COL[7929] = 1'b0;
assign COL[7930] = 1'b1;
assign COL[7931] = 1'b1;
assign COL[7932] = 1'b1;
assign COL[7933] = 1'b1;
assign COL[7934] = 1'b1;
assign COL[7935] = 1'b0;
assign COL[7936] = 1'b0;
assign COL[7937] = 1'b0;
assign COL[7938] = 1'b0;
assign COL[7939] = 1'b0;
assign COL[7940] = 1'b0;
assign COL[7941] = 1'b0;
assign COL[7942] = 1'b0;
assign COL[7943] = 1'b0;
assign COL[7944] = 1'b0;
assign COL[7945] = 1'b0;
assign COL[7946] = 1'b0;
assign COL[7947] = 1'b0;
assign COL[7948] = 1'b0;
assign COL[7949] = 1'b0;
assign COL[7950] = 1'b0;
assign COL[7951] = 1'b0;
assign COL[7952] = 1'b0;
assign COL[7953] = 1'b0;
assign COL[7954] = 1'b0;
assign COL[7955] = 1'b0;
assign COL[7956] = 1'b0;
assign COL[7957] = 1'b0;
assign COL[7958] = 1'b0;
assign COL[7959] = 1'b0;
assign COL[7960] = 1'b0;
assign COL[7961] = 1'b0;
assign COL[7962] = 1'b0;
assign COL[7963] = 1'b0;
assign COL[7964] = 1'b0;
assign COL[7965] = 1'b0;
assign COL[7966] = 1'b0;
assign COL[7967] = 1'b0;
assign COL[7968] = 1'b0;
assign COL[7969] = 1'b0;
assign COL[7970] = 1'b0;
assign COL[7971] = 1'b0;
assign COL[7972] = 1'b0;
assign COL[7973] = 1'b0;
assign COL[7974] = 1'b0;
assign COL[7975] = 1'b0;
assign COL[7976] = 1'b0;
assign COL[7977] = 1'b0;
assign COL[7978] = 1'b0;
assign COL[7979] = 1'b0;
assign COL[7980] = 1'b0;
assign COL[7981] = 1'b0;
assign COL[7982] = 1'b0;
assign COL[7983] = 1'b0;
assign COL[7984] = 1'b0;
assign COL[7985] = 1'b0;
assign COL[7986] = 1'b0;
assign COL[7987] = 1'b0;
assign COL[7988] = 1'b0;
assign COL[7989] = 1'b0;
assign COL[7990] = 1'b0;
assign COL[7991] = 1'b0;
assign COL[7992] = 1'b0;
assign COL[7993] = 1'b0;
assign COL[7994] = 1'b0;
assign COL[7995] = 1'b0;
assign COL[7996] = 1'b0;
assign COL[7997] = 1'b0;
assign COL[7998] = 1'b0;
assign COL[7999] = 1'b0;
assign COL[8000] = 1'b0;
assign COL[8001] = 1'b1;
assign COL[8002] = 1'b1;
assign COL[8003] = 1'b1;
assign COL[8004] = 1'b1;
assign COL[8005] = 1'b1;
assign COL[8006] = 1'b0;
assign COL[8007] = 1'b0;
assign COL[8008] = 1'b0;
assign COL[8009] = 1'b0;
assign COL[8010] = 1'b0;
assign COL[8011] = 1'b0;
assign COL[8012] = 1'b0;
assign COL[8013] = 1'b0;
assign COL[8014] = 1'b0;
assign COL[8015] = 1'b0;
assign COL[8016] = 1'b1;
assign COL[8017] = 1'b1;
assign COL[8018] = 1'b1;
assign COL[8019] = 1'b1;
assign COL[8020] = 1'b1;
assign COL[8021] = 1'b1;
assign COL[8022] = 1'b1;
assign COL[8023] = 1'b1;
assign COL[8024] = 1'b1;
assign COL[8025] = 1'b1;
assign COL[8026] = 1'b1;
assign COL[8027] = 1'b1;
assign COL[8028] = 1'b1;
assign COL[8029] = 1'b1;
assign COL[8030] = 1'b1;
assign COL[8031] = 1'b1;
assign COL[8032] = 1'b1;
assign COL[8033] = 1'b1;
assign COL[8034] = 1'b1;
assign COL[8035] = 1'b1;
assign COL[8036] = 1'b1;
assign COL[8037] = 1'b1;
assign COL[8038] = 1'b1;
assign COL[8039] = 1'b1;
assign COL[8040] = 1'b1;
assign COL[8041] = 1'b1;
assign COL[8042] = 1'b1;
assign COL[8043] = 1'b1;
assign COL[8044] = 1'b1;
assign COL[8045] = 1'b1;
assign COL[8046] = 1'b1;
assign COL[8047] = 1'b1;
assign COL[8048] = 1'b1;
assign COL[8049] = 1'b1;
assign COL[8050] = 1'b1;
assign COL[8051] = 1'b1;
assign COL[8052] = 1'b1;
assign COL[8053] = 1'b1;
assign COL[8054] = 1'b1;
assign COL[8055] = 1'b1;
assign COL[8056] = 1'b1;
assign COL[8057] = 1'b1;
assign COL[8058] = 1'b1;
assign COL[8059] = 1'b1;
assign COL[8060] = 1'b1;
assign COL[8061] = 1'b1;
assign COL[8062] = 1'b0;
assign COL[8063] = 1'b0;
assign COL[8064] = 1'b0;
assign COL[8065] = 1'b0;
assign COL[8066] = 1'b0;
assign COL[8067] = 1'b0;
assign COL[8068] = 1'b0;
assign COL[8069] = 1'b0;
assign COL[8070] = 1'b1;
assign COL[8071] = 1'b1;
assign COL[8072] = 1'b1;
assign COL[8073] = 1'b1;
assign COL[8074] = 1'b1;
assign COL[8075] = 1'b0;
assign COL[8076] = 1'b0;
assign COL[8077] = 1'b0;
assign COL[8078] = 1'b0;
assign COL[8079] = 1'b0;
assign COL[8080] = 1'b0;
assign COL[8081] = 1'b0;
assign COL[8082] = 1'b0;
assign COL[8083] = 1'b0;
assign COL[8084] = 1'b0;
assign COL[8085] = 1'b0;
assign COL[8086] = 1'b0;
assign COL[8087] = 1'b0;
assign COL[8088] = 1'b0;
assign COL[8089] = 1'b0;
assign COL[8090] = 1'b1;
assign COL[8091] = 1'b1;
assign COL[8092] = 1'b1;
assign COL[8093] = 1'b1;
assign COL[8094] = 1'b1;
assign COL[8095] = 1'b0;
assign COL[8096] = 1'b0;
assign COL[8097] = 1'b0;
assign COL[8098] = 1'b0;
assign COL[8099] = 1'b0;
assign COL[8100] = 1'b0;
assign COL[8101] = 1'b0;
assign COL[8102] = 1'b0;
assign COL[8103] = 1'b0;
assign COL[8104] = 1'b0;
assign COL[8105] = 1'b0;
assign COL[8106] = 1'b0;
assign COL[8107] = 1'b0;
assign COL[8108] = 1'b0;
assign COL[8109] = 1'b0;
assign COL[8110] = 1'b0;
assign COL[8111] = 1'b0;
assign COL[8112] = 1'b0;
assign COL[8113] = 1'b0;
assign COL[8114] = 1'b0;
assign COL[8115] = 1'b0;
assign COL[8116] = 1'b0;
assign COL[8117] = 1'b0;
assign COL[8118] = 1'b0;
assign COL[8119] = 1'b0;
assign COL[8120] = 1'b0;
assign COL[8121] = 1'b0;
assign COL[8122] = 1'b0;
assign COL[8123] = 1'b0;
assign COL[8124] = 1'b0;
assign COL[8125] = 1'b0;
assign COL[8126] = 1'b0;
assign COL[8127] = 1'b0;
assign COL[8128] = 1'b0;
assign COL[8129] = 1'b0;
assign COL[8130] = 1'b0;
assign COL[8131] = 1'b0;
assign COL[8132] = 1'b0;
assign COL[8133] = 1'b0;
assign COL[8134] = 1'b0;
assign COL[8135] = 1'b0;
assign COL[8136] = 1'b0;
assign COL[8137] = 1'b0;
assign COL[8138] = 1'b0;
assign COL[8139] = 1'b0;
assign COL[8140] = 1'b0;
assign COL[8141] = 1'b0;
assign COL[8142] = 1'b0;
assign COL[8143] = 1'b0;
assign COL[8144] = 1'b0;
assign COL[8145] = 1'b0;
assign COL[8146] = 1'b0;
assign COL[8147] = 1'b0;
assign COL[8148] = 1'b0;
assign COL[8149] = 1'b0;
assign COL[8150] = 1'b0;
assign COL[8151] = 1'b0;
assign COL[8152] = 1'b0;
assign COL[8153] = 1'b0;
assign COL[8154] = 1'b0;
assign COL[8155] = 1'b0;
assign COL[8156] = 1'b0;
assign COL[8157] = 1'b0;
assign COL[8158] = 1'b0;
assign COL[8159] = 1'b0;
assign COL[8160] = 1'b0;
assign COL[8161] = 1'b1;
assign COL[8162] = 1'b1;
assign COL[8163] = 1'b1;
assign COL[8164] = 1'b1;
assign COL[8165] = 1'b1;
assign COL[8166] = 1'b0;
assign COL[8167] = 1'b0;
assign COL[8168] = 1'b0;
assign COL[8169] = 1'b0;
assign COL[8170] = 1'b0;
assign COL[8171] = 1'b0;
assign COL[8172] = 1'b0;
assign COL[8173] = 1'b0;
assign COL[8174] = 1'b0;
assign COL[8175] = 1'b0;
assign COL[8176] = 1'b0;
assign COL[8177] = 1'b0;
assign COL[8178] = 1'b0;
assign COL[8179] = 1'b0;
assign COL[8180] = 1'b0;
assign COL[8181] = 1'b0;
assign COL[8182] = 1'b0;
assign COL[8183] = 1'b0;
assign COL[8184] = 1'b0;
assign COL[8185] = 1'b0;
assign COL[8186] = 1'b0;
assign COL[8187] = 1'b0;
assign COL[8188] = 1'b0;
assign COL[8189] = 1'b1;
assign COL[8190] = 1'b1;
assign COL[8191] = 1'b1;
assign COL[8192] = 1'b1;
assign COL[8193] = 1'b0;
assign COL[8194] = 1'b0;
assign COL[8195] = 1'b0;
assign COL[8196] = 1'b0;
assign COL[8197] = 1'b0;
assign COL[8198] = 1'b0;
assign COL[8199] = 1'b0;
assign COL[8200] = 1'b0;
assign COL[8201] = 1'b0;
assign COL[8202] = 1'b0;
assign COL[8203] = 1'b0;
assign COL[8204] = 1'b0;
assign COL[8205] = 1'b0;
assign COL[8206] = 1'b0;
assign COL[8207] = 1'b0;
assign COL[8208] = 1'b0;
assign COL[8209] = 1'b0;
assign COL[8210] = 1'b0;
assign COL[8211] = 1'b0;
assign COL[8212] = 1'b0;
assign COL[8213] = 1'b0;
assign COL[8214] = 1'b0;
assign COL[8215] = 1'b0;
assign COL[8216] = 1'b0;
assign COL[8217] = 1'b0;
assign COL[8218] = 1'b1;
assign COL[8219] = 1'b1;
assign COL[8220] = 1'b1;
assign COL[8221] = 1'b1;
assign COL[8222] = 1'b0;
assign COL[8223] = 1'b0;
assign COL[8224] = 1'b0;
assign COL[8225] = 1'b0;
assign COL[8226] = 1'b0;
assign COL[8227] = 1'b0;
assign COL[8228] = 1'b0;
assign COL[8229] = 1'b0;
assign COL[8230] = 1'b1;
assign COL[8231] = 1'b1;
assign COL[8232] = 1'b1;
assign COL[8233] = 1'b1;
assign COL[8234] = 1'b1;
assign COL[8235] = 1'b0;
assign COL[8236] = 1'b0;
assign COL[8237] = 1'b0;
assign COL[8238] = 1'b0;
assign COL[8239] = 1'b0;
assign COL[8240] = 1'b0;
assign COL[8241] = 1'b0;
assign COL[8242] = 1'b0;
assign COL[8243] = 1'b0;
assign COL[8244] = 1'b0;
assign COL[8245] = 1'b0;
assign COL[8246] = 1'b0;
assign COL[8247] = 1'b0;
assign COL[8248] = 1'b0;
assign COL[8249] = 1'b0;
assign COL[8250] = 1'b1;
assign COL[8251] = 1'b1;
assign COL[8252] = 1'b1;
assign COL[8253] = 1'b1;
assign COL[8254] = 1'b1;
assign COL[8255] = 1'b0;
assign COL[8256] = 1'b0;
assign COL[8257] = 1'b0;
assign COL[8258] = 1'b0;
assign COL[8259] = 1'b0;
assign COL[8260] = 1'b0;
assign COL[8261] = 1'b0;
assign COL[8262] = 1'b0;
assign COL[8263] = 1'b0;
assign COL[8264] = 1'b0;
assign COL[8265] = 1'b0;
assign COL[8266] = 1'b0;
assign COL[8267] = 1'b0;
assign COL[8268] = 1'b0;
assign COL[8269] = 1'b0;
assign COL[8270] = 1'b0;
assign COL[8271] = 1'b0;
assign COL[8272] = 1'b0;
assign COL[8273] = 1'b0;
assign COL[8274] = 1'b0;
assign COL[8275] = 1'b0;
assign COL[8276] = 1'b0;
assign COL[8277] = 1'b0;
assign COL[8278] = 1'b0;
assign COL[8279] = 1'b0;
assign COL[8280] = 1'b0;
assign COL[8281] = 1'b0;
assign COL[8282] = 1'b0;
assign COL[8283] = 1'b0;
assign COL[8284] = 1'b0;
assign COL[8285] = 1'b0;
assign COL[8286] = 1'b0;
assign COL[8287] = 1'b0;
assign COL[8288] = 1'b0;
assign COL[8289] = 1'b0;
assign COL[8290] = 1'b0;
assign COL[8291] = 1'b0;
assign COL[8292] = 1'b0;
assign COL[8293] = 1'b0;
assign COL[8294] = 1'b0;
assign COL[8295] = 1'b0;
assign COL[8296] = 1'b0;
assign COL[8297] = 1'b0;
assign COL[8298] = 1'b0;
assign COL[8299] = 1'b0;
assign COL[8300] = 1'b0;
assign COL[8301] = 1'b0;
assign COL[8302] = 1'b0;
assign COL[8303] = 1'b0;
assign COL[8304] = 1'b0;
assign COL[8305] = 1'b0;
assign COL[8306] = 1'b0;
assign COL[8307] = 1'b0;
assign COL[8308] = 1'b0;
assign COL[8309] = 1'b0;
assign COL[8310] = 1'b0;
assign COL[8311] = 1'b0;
assign COL[8312] = 1'b0;
assign COL[8313] = 1'b0;
assign COL[8314] = 1'b0;
assign COL[8315] = 1'b0;
assign COL[8316] = 1'b0;
assign COL[8317] = 1'b0;
assign COL[8318] = 1'b0;
assign COL[8319] = 1'b0;
assign COL[8320] = 1'b0;
assign COL[8321] = 1'b1;
assign COL[8322] = 1'b1;
assign COL[8323] = 1'b1;
assign COL[8324] = 1'b1;
assign COL[8325] = 1'b1;
assign COL[8326] = 1'b0;
assign COL[8327] = 1'b0;
assign COL[8328] = 1'b0;
assign COL[8329] = 1'b0;
assign COL[8330] = 1'b0;
assign COL[8331] = 1'b0;
assign COL[8332] = 1'b0;
assign COL[8333] = 1'b0;
assign COL[8334] = 1'b0;
assign COL[8335] = 1'b0;
assign COL[8336] = 1'b0;
assign COL[8337] = 1'b0;
assign COL[8338] = 1'b0;
assign COL[8339] = 1'b0;
assign COL[8340] = 1'b0;
assign COL[8341] = 1'b0;
assign COL[8342] = 1'b0;
assign COL[8343] = 1'b0;
assign COL[8344] = 1'b0;
assign COL[8345] = 1'b0;
assign COL[8346] = 1'b0;
assign COL[8347] = 1'b0;
assign COL[8348] = 1'b0;
assign COL[8349] = 1'b1;
assign COL[8350] = 1'b1;
assign COL[8351] = 1'b1;
assign COL[8352] = 1'b1;
assign COL[8353] = 1'b0;
assign COL[8354] = 1'b0;
assign COL[8355] = 1'b0;
assign COL[8356] = 1'b0;
assign COL[8357] = 1'b0;
assign COL[8358] = 1'b0;
assign COL[8359] = 1'b0;
assign COL[8360] = 1'b0;
assign COL[8361] = 1'b0;
assign COL[8362] = 1'b0;
assign COL[8363] = 1'b0;
assign COL[8364] = 1'b0;
assign COL[8365] = 1'b0;
assign COL[8366] = 1'b0;
assign COL[8367] = 1'b0;
assign COL[8368] = 1'b0;
assign COL[8369] = 1'b0;
assign COL[8370] = 1'b0;
assign COL[8371] = 1'b0;
assign COL[8372] = 1'b0;
assign COL[8373] = 1'b0;
assign COL[8374] = 1'b0;
assign COL[8375] = 1'b0;
assign COL[8376] = 1'b0;
assign COL[8377] = 1'b0;
assign COL[8378] = 1'b1;
assign COL[8379] = 1'b1;
assign COL[8380] = 1'b1;
assign COL[8381] = 1'b1;
assign COL[8382] = 1'b0;
assign COL[8383] = 1'b0;
assign COL[8384] = 1'b0;
assign COL[8385] = 1'b0;
assign COL[8386] = 1'b0;
assign COL[8387] = 1'b0;
assign COL[8388] = 1'b0;
assign COL[8389] = 1'b0;
assign COL[8390] = 1'b1;
assign COL[8391] = 1'b1;
assign COL[8392] = 1'b1;
assign COL[8393] = 1'b1;
assign COL[8394] = 1'b1;
assign COL[8395] = 1'b0;
assign COL[8396] = 1'b0;
assign COL[8397] = 1'b0;
assign COL[8398] = 1'b0;
assign COL[8399] = 1'b0;
assign COL[8400] = 1'b0;
assign COL[8401] = 1'b0;
assign COL[8402] = 1'b0;
assign COL[8403] = 1'b0;
assign COL[8404] = 1'b0;
assign COL[8405] = 1'b0;
assign COL[8406] = 1'b0;
assign COL[8407] = 1'b0;
assign COL[8408] = 1'b0;
assign COL[8409] = 1'b0;
assign COL[8410] = 1'b1;
assign COL[8411] = 1'b1;
assign COL[8412] = 1'b1;
assign COL[8413] = 1'b1;
assign COL[8414] = 1'b1;
assign COL[8415] = 1'b0;
assign COL[8416] = 1'b0;
assign COL[8417] = 1'b0;
assign COL[8418] = 1'b0;
assign COL[8419] = 1'b0;
assign COL[8420] = 1'b0;
assign COL[8421] = 1'b0;
assign COL[8422] = 1'b0;
assign COL[8423] = 1'b0;
assign COL[8424] = 1'b0;
assign COL[8425] = 1'b0;
assign COL[8426] = 1'b0;
assign COL[8427] = 1'b0;
assign COL[8428] = 1'b0;
assign COL[8429] = 1'b0;
assign COL[8430] = 1'b0;
assign COL[8431] = 1'b0;
assign COL[8432] = 1'b0;
assign COL[8433] = 1'b0;
assign COL[8434] = 1'b0;
assign COL[8435] = 1'b0;
assign COL[8436] = 1'b0;
assign COL[8437] = 1'b0;
assign COL[8438] = 1'b0;
assign COL[8439] = 1'b0;
assign COL[8440] = 1'b0;
assign COL[8441] = 1'b0;
assign COL[8442] = 1'b0;
assign COL[8443] = 1'b0;
assign COL[8444] = 1'b0;
assign COL[8445] = 1'b0;
assign COL[8446] = 1'b0;
assign COL[8447] = 1'b0;
assign COL[8448] = 1'b0;
assign COL[8449] = 1'b0;
assign COL[8450] = 1'b0;
assign COL[8451] = 1'b0;
assign COL[8452] = 1'b0;
assign COL[8453] = 1'b0;
assign COL[8454] = 1'b0;
assign COL[8455] = 1'b0;
assign COL[8456] = 1'b0;
assign COL[8457] = 1'b0;
assign COL[8458] = 1'b0;
assign COL[8459] = 1'b0;
assign COL[8460] = 1'b0;
assign COL[8461] = 1'b0;
assign COL[8462] = 1'b0;
assign COL[8463] = 1'b0;
assign COL[8464] = 1'b0;
assign COL[8465] = 1'b0;
assign COL[8466] = 1'b0;
assign COL[8467] = 1'b0;
assign COL[8468] = 1'b0;
assign COL[8469] = 1'b0;
assign COL[8470] = 1'b0;
assign COL[8471] = 1'b0;
assign COL[8472] = 1'b0;
assign COL[8473] = 1'b0;
assign COL[8474] = 1'b0;
assign COL[8475] = 1'b0;
assign COL[8476] = 1'b0;
assign COL[8477] = 1'b0;
assign COL[8478] = 1'b0;
assign COL[8479] = 1'b0;
assign COL[8480] = 1'b0;
assign COL[8481] = 1'b1;
assign COL[8482] = 1'b1;
assign COL[8483] = 1'b1;
assign COL[8484] = 1'b1;
assign COL[8485] = 1'b1;
assign COL[8486] = 1'b0;
assign COL[8487] = 1'b0;
assign COL[8488] = 1'b0;
assign COL[8489] = 1'b0;
assign COL[8490] = 1'b0;
assign COL[8491] = 1'b0;
assign COL[8492] = 1'b0;
assign COL[8493] = 1'b0;
assign COL[8494] = 1'b0;
assign COL[8495] = 1'b0;
assign COL[8496] = 1'b0;
assign COL[8497] = 1'b0;
assign COL[8498] = 1'b0;
assign COL[8499] = 1'b0;
assign COL[8500] = 1'b0;
assign COL[8501] = 1'b0;
assign COL[8502] = 1'b0;
assign COL[8503] = 1'b0;
assign COL[8504] = 1'b0;
assign COL[8505] = 1'b0;
assign COL[8506] = 1'b0;
assign COL[8507] = 1'b0;
assign COL[8508] = 1'b0;
assign COL[8509] = 1'b1;
assign COL[8510] = 1'b1;
assign COL[8511] = 1'b1;
assign COL[8512] = 1'b1;
assign COL[8513] = 1'b0;
assign COL[8514] = 1'b0;
assign COL[8515] = 1'b0;
assign COL[8516] = 1'b0;
assign COL[8517] = 1'b0;
assign COL[8518] = 1'b0;
assign COL[8519] = 1'b0;
assign COL[8520] = 1'b0;
assign COL[8521] = 1'b0;
assign COL[8522] = 1'b0;
assign COL[8523] = 1'b0;
assign COL[8524] = 1'b0;
assign COL[8525] = 1'b0;
assign COL[8526] = 1'b0;
assign COL[8527] = 1'b0;
assign COL[8528] = 1'b0;
assign COL[8529] = 1'b0;
assign COL[8530] = 1'b0;
assign COL[8531] = 1'b0;
assign COL[8532] = 1'b0;
assign COL[8533] = 1'b0;
assign COL[8534] = 1'b0;
assign COL[8535] = 1'b0;
assign COL[8536] = 1'b0;
assign COL[8537] = 1'b0;
assign COL[8538] = 1'b1;
assign COL[8539] = 1'b1;
assign COL[8540] = 1'b1;
assign COL[8541] = 1'b1;
assign COL[8542] = 1'b0;
assign COL[8543] = 1'b0;
assign COL[8544] = 1'b0;
assign COL[8545] = 1'b0;
assign COL[8546] = 1'b0;
assign COL[8547] = 1'b0;
assign COL[8548] = 1'b0;
assign COL[8549] = 1'b0;
assign COL[8550] = 1'b1;
assign COL[8551] = 1'b1;
assign COL[8552] = 1'b1;
assign COL[8553] = 1'b1;
assign COL[8554] = 1'b1;
assign COL[8555] = 1'b0;
assign COL[8556] = 1'b0;
assign COL[8557] = 1'b0;
assign COL[8558] = 1'b0;
assign COL[8559] = 1'b0;
assign COL[8560] = 1'b0;
assign COL[8561] = 1'b0;
assign COL[8562] = 1'b0;
assign COL[8563] = 1'b0;
assign COL[8564] = 1'b0;
assign COL[8565] = 1'b0;
assign COL[8566] = 1'b0;
assign COL[8567] = 1'b0;
assign COL[8568] = 1'b0;
assign COL[8569] = 1'b0;
assign COL[8570] = 1'b1;
assign COL[8571] = 1'b1;
assign COL[8572] = 1'b1;
assign COL[8573] = 1'b1;
assign COL[8574] = 1'b1;
assign COL[8575] = 1'b0;
assign COL[8576] = 1'b0;
assign COL[8577] = 1'b0;
assign COL[8578] = 1'b0;
assign COL[8579] = 1'b0;
assign COL[8580] = 1'b0;
assign COL[8581] = 1'b0;
assign COL[8582] = 1'b0;
assign COL[8583] = 1'b0;
assign COL[8584] = 1'b0;
assign COL[8585] = 1'b0;
assign COL[8586] = 1'b0;
assign COL[8587] = 1'b0;
assign COL[8588] = 1'b0;
assign COL[8589] = 1'b0;
assign COL[8590] = 1'b0;
assign COL[8591] = 1'b0;
assign COL[8592] = 1'b0;
assign COL[8593] = 1'b0;
assign COL[8594] = 1'b0;
assign COL[8595] = 1'b0;
assign COL[8596] = 1'b0;
assign COL[8597] = 1'b0;
assign COL[8598] = 1'b0;
assign COL[8599] = 1'b0;
assign COL[8600] = 1'b0;
assign COL[8601] = 1'b0;
assign COL[8602] = 1'b0;
assign COL[8603] = 1'b0;
assign COL[8604] = 1'b0;
assign COL[8605] = 1'b0;
assign COL[8606] = 1'b0;
assign COL[8607] = 1'b0;
assign COL[8608] = 1'b0;
assign COL[8609] = 1'b0;
assign COL[8610] = 1'b0;
assign COL[8611] = 1'b0;
assign COL[8612] = 1'b0;
assign COL[8613] = 1'b0;
assign COL[8614] = 1'b0;
assign COL[8615] = 1'b0;
assign COL[8616] = 1'b0;
assign COL[8617] = 1'b0;
assign COL[8618] = 1'b0;
assign COL[8619] = 1'b0;
assign COL[8620] = 1'b0;
assign COL[8621] = 1'b0;
assign COL[8622] = 1'b0;
assign COL[8623] = 1'b0;
assign COL[8624] = 1'b0;
assign COL[8625] = 1'b0;
assign COL[8626] = 1'b0;
assign COL[8627] = 1'b0;
assign COL[8628] = 1'b0;
assign COL[8629] = 1'b0;
assign COL[8630] = 1'b0;
assign COL[8631] = 1'b0;
assign COL[8632] = 1'b0;
assign COL[8633] = 1'b0;
assign COL[8634] = 1'b0;
assign COL[8635] = 1'b0;
assign COL[8636] = 1'b0;
assign COL[8637] = 1'b0;
assign COL[8638] = 1'b0;
assign COL[8639] = 1'b0;
assign COL[8640] = 1'b0;
assign COL[8641] = 1'b1;
assign COL[8642] = 1'b1;
assign COL[8643] = 1'b1;
assign COL[8644] = 1'b1;
assign COL[8645] = 1'b1;
assign COL[8646] = 1'b0;
assign COL[8647] = 1'b0;
assign COL[8648] = 1'b0;
assign COL[8649] = 1'b0;
assign COL[8650] = 1'b0;
assign COL[8651] = 1'b0;
assign COL[8652] = 1'b0;
assign COL[8653] = 1'b0;
assign COL[8654] = 1'b0;
assign COL[8655] = 1'b0;
assign COL[8656] = 1'b0;
assign COL[8657] = 1'b0;
assign COL[8658] = 1'b0;
assign COL[8659] = 1'b0;
assign COL[8660] = 1'b0;
assign COL[8661] = 1'b0;
assign COL[8662] = 1'b0;
assign COL[8663] = 1'b0;
assign COL[8664] = 1'b0;
assign COL[8665] = 1'b0;
assign COL[8666] = 1'b0;
assign COL[8667] = 1'b0;
assign COL[8668] = 1'b0;
assign COL[8669] = 1'b1;
assign COL[8670] = 1'b1;
assign COL[8671] = 1'b1;
assign COL[8672] = 1'b1;
assign COL[8673] = 1'b0;
assign COL[8674] = 1'b0;
assign COL[8675] = 1'b0;
assign COL[8676] = 1'b0;
assign COL[8677] = 1'b0;
assign COL[8678] = 1'b0;
assign COL[8679] = 1'b0;
assign COL[8680] = 1'b0;
assign COL[8681] = 1'b0;
assign COL[8682] = 1'b0;
assign COL[8683] = 1'b0;
assign COL[8684] = 1'b0;
assign COL[8685] = 1'b0;
assign COL[8686] = 1'b0;
assign COL[8687] = 1'b0;
assign COL[8688] = 1'b0;
assign COL[8689] = 1'b0;
assign COL[8690] = 1'b0;
assign COL[8691] = 1'b0;
assign COL[8692] = 1'b0;
assign COL[8693] = 1'b0;
assign COL[8694] = 1'b0;
assign COL[8695] = 1'b0;
assign COL[8696] = 1'b0;
assign COL[8697] = 1'b0;
assign COL[8698] = 1'b1;
assign COL[8699] = 1'b1;
assign COL[8700] = 1'b1;
assign COL[8701] = 1'b1;
assign COL[8702] = 1'b0;
assign COL[8703] = 1'b0;
assign COL[8704] = 1'b0;
assign COL[8705] = 1'b0;
assign COL[8706] = 1'b0;
assign COL[8707] = 1'b0;
assign COL[8708] = 1'b0;
assign COL[8709] = 1'b0;
assign COL[8710] = 1'b1;
assign COL[8711] = 1'b1;
assign COL[8712] = 1'b1;
assign COL[8713] = 1'b1;
assign COL[8714] = 1'b1;
assign COL[8715] = 1'b0;
assign COL[8716] = 1'b0;
assign COL[8717] = 1'b0;
assign COL[8718] = 1'b0;
assign COL[8719] = 1'b0;
assign COL[8720] = 1'b0;
assign COL[8721] = 1'b0;
assign COL[8722] = 1'b0;
assign COL[8723] = 1'b0;
assign COL[8724] = 1'b0;
assign COL[8725] = 1'b0;
assign COL[8726] = 1'b0;
assign COL[8727] = 1'b0;
assign COL[8728] = 1'b0;
assign COL[8729] = 1'b0;
assign COL[8730] = 1'b1;
assign COL[8731] = 1'b1;
assign COL[8732] = 1'b1;
assign COL[8733] = 1'b1;
assign COL[8734] = 1'b1;
assign COL[8735] = 1'b0;
assign COL[8736] = 1'b0;
assign COL[8737] = 1'b0;
assign COL[8738] = 1'b0;
assign COL[8739] = 1'b0;
assign COL[8740] = 1'b0;
assign COL[8741] = 1'b0;
assign COL[8742] = 1'b0;
assign COL[8743] = 1'b0;
assign COL[8744] = 1'b0;
assign COL[8745] = 1'b0;
assign COL[8746] = 1'b0;
assign COL[8747] = 1'b0;
assign COL[8748] = 1'b0;
assign COL[8749] = 1'b0;
assign COL[8750] = 1'b0;
assign COL[8751] = 1'b0;
assign COL[8752] = 1'b0;
assign COL[8753] = 1'b0;
assign COL[8754] = 1'b0;
assign COL[8755] = 1'b0;
assign COL[8756] = 1'b0;
assign COL[8757] = 1'b0;
assign COL[8758] = 1'b0;
assign COL[8759] = 1'b0;
assign COL[8760] = 1'b0;
assign COL[8761] = 1'b0;
assign COL[8762] = 1'b0;
assign COL[8763] = 1'b0;
assign COL[8764] = 1'b0;
assign COL[8765] = 1'b0;
assign COL[8766] = 1'b0;
assign COL[8767] = 1'b0;
assign COL[8768] = 1'b0;
assign COL[8769] = 1'b0;
assign COL[8770] = 1'b0;
assign COL[8771] = 1'b0;
assign COL[8772] = 1'b0;
assign COL[8773] = 1'b0;
assign COL[8774] = 1'b0;
assign COL[8775] = 1'b0;
assign COL[8776] = 1'b0;
assign COL[8777] = 1'b0;
assign COL[8778] = 1'b0;
assign COL[8779] = 1'b0;
assign COL[8780] = 1'b0;
assign COL[8781] = 1'b0;
assign COL[8782] = 1'b0;
assign COL[8783] = 1'b0;
assign COL[8784] = 1'b0;
assign COL[8785] = 1'b0;
assign COL[8786] = 1'b0;
assign COL[8787] = 1'b0;
assign COL[8788] = 1'b0;
assign COL[8789] = 1'b0;
assign COL[8790] = 1'b0;
assign COL[8791] = 1'b0;
assign COL[8792] = 1'b0;
assign COL[8793] = 1'b0;
assign COL[8794] = 1'b0;
assign COL[8795] = 1'b0;
assign COL[8796] = 1'b0;
assign COL[8797] = 1'b0;
assign COL[8798] = 1'b0;
assign COL[8799] = 1'b0;
assign COL[8800] = 1'b0;
assign COL[8801] = 1'b1;
assign COL[8802] = 1'b1;
assign COL[8803] = 1'b1;
assign COL[8804] = 1'b1;
assign COL[8805] = 1'b1;
assign COL[8806] = 1'b0;
assign COL[8807] = 1'b0;
assign COL[8808] = 1'b0;
assign COL[8809] = 1'b0;
assign COL[8810] = 1'b0;
assign COL[8811] = 1'b0;
assign COL[8812] = 1'b0;
assign COL[8813] = 1'b0;
assign COL[8814] = 1'b0;
assign COL[8815] = 1'b0;
assign COL[8816] = 1'b0;
assign COL[8817] = 1'b0;
assign COL[8818] = 1'b0;
assign COL[8819] = 1'b0;
assign COL[8820] = 1'b0;
assign COL[8821] = 1'b0;
assign COL[8822] = 1'b0;
assign COL[8823] = 1'b0;
assign COL[8824] = 1'b0;
assign COL[8825] = 1'b0;
assign COL[8826] = 1'b0;
assign COL[8827] = 1'b0;
assign COL[8828] = 1'b0;
assign COL[8829] = 1'b1;
assign COL[8830] = 1'b1;
assign COL[8831] = 1'b1;
assign COL[8832] = 1'b1;
assign COL[8833] = 1'b0;
assign COL[8834] = 1'b0;
assign COL[8835] = 1'b0;
assign COL[8836] = 1'b0;
assign COL[8837] = 1'b0;
assign COL[8838] = 1'b0;
assign COL[8839] = 1'b0;
assign COL[8840] = 1'b0;
assign COL[8841] = 1'b0;
assign COL[8842] = 1'b0;
assign COL[8843] = 1'b0;
assign COL[8844] = 1'b0;
assign COL[8845] = 1'b0;
assign COL[8846] = 1'b0;
assign COL[8847] = 1'b0;
assign COL[8848] = 1'b0;
assign COL[8849] = 1'b0;
assign COL[8850] = 1'b0;
assign COL[8851] = 1'b0;
assign COL[8852] = 1'b0;
assign COL[8853] = 1'b0;
assign COL[8854] = 1'b0;
assign COL[8855] = 1'b0;
assign COL[8856] = 1'b0;
assign COL[8857] = 1'b0;
assign COL[8858] = 1'b1;
assign COL[8859] = 1'b1;
assign COL[8860] = 1'b1;
assign COL[8861] = 1'b1;
assign COL[8862] = 1'b0;
assign COL[8863] = 1'b0;
assign COL[8864] = 1'b0;
assign COL[8865] = 1'b0;
assign COL[8866] = 1'b0;
assign COL[8867] = 1'b0;
assign COL[8868] = 1'b0;
assign COL[8869] = 1'b0;
assign COL[8870] = 1'b1;
assign COL[8871] = 1'b1;
assign COL[8872] = 1'b1;
assign COL[8873] = 1'b1;
assign COL[8874] = 1'b1;
assign COL[8875] = 1'b0;
assign COL[8876] = 1'b0;
assign COL[8877] = 1'b0;
assign COL[8878] = 1'b0;
assign COL[8879] = 1'b0;
assign COL[8880] = 1'b0;
assign COL[8881] = 1'b0;
assign COL[8882] = 1'b0;
assign COL[8883] = 1'b0;
assign COL[8884] = 1'b0;
assign COL[8885] = 1'b0;
assign COL[8886] = 1'b0;
assign COL[8887] = 1'b0;
assign COL[8888] = 1'b0;
assign COL[8889] = 1'b0;
assign COL[8890] = 1'b1;
assign COL[8891] = 1'b1;
assign COL[8892] = 1'b1;
assign COL[8893] = 1'b1;
assign COL[8894] = 1'b1;
assign COL[8895] = 1'b0;
assign COL[8896] = 1'b0;
assign COL[8897] = 1'b0;
assign COL[8898] = 1'b0;
assign COL[8899] = 1'b0;
assign COL[8900] = 1'b0;
assign COL[8901] = 1'b0;
assign COL[8902] = 1'b0;
assign COL[8903] = 1'b0;
assign COL[8904] = 1'b0;
assign COL[8905] = 1'b0;
assign COL[8906] = 1'b0;
assign COL[8907] = 1'b0;
assign COL[8908] = 1'b0;
assign COL[8909] = 1'b0;
assign COL[8910] = 1'b0;
assign COL[8911] = 1'b0;
assign COL[8912] = 1'b0;
assign COL[8913] = 1'b0;
assign COL[8914] = 1'b0;
assign COL[8915] = 1'b0;
assign COL[8916] = 1'b0;
assign COL[8917] = 1'b0;
assign COL[8918] = 1'b0;
assign COL[8919] = 1'b0;
assign COL[8920] = 1'b0;
assign COL[8921] = 1'b0;
assign COL[8922] = 1'b0;
assign COL[8923] = 1'b0;
assign COL[8924] = 1'b0;
assign COL[8925] = 1'b0;
assign COL[8926] = 1'b0;
assign COL[8927] = 1'b0;
assign COL[8928] = 1'b0;
assign COL[8929] = 1'b0;
assign COL[8930] = 1'b0;
assign COL[8931] = 1'b0;
assign COL[8932] = 1'b0;
assign COL[8933] = 1'b0;
assign COL[8934] = 1'b0;
assign COL[8935] = 1'b0;
assign COL[8936] = 1'b0;
assign COL[8937] = 1'b0;
assign COL[8938] = 1'b0;
assign COL[8939] = 1'b0;
assign COL[8940] = 1'b0;
assign COL[8941] = 1'b0;
assign COL[8942] = 1'b0;
assign COL[8943] = 1'b0;
assign COL[8944] = 1'b0;
assign COL[8945] = 1'b0;
assign COL[8946] = 1'b0;
assign COL[8947] = 1'b0;
assign COL[8948] = 1'b0;
assign COL[8949] = 1'b0;
assign COL[8950] = 1'b0;
assign COL[8951] = 1'b0;
assign COL[8952] = 1'b0;
assign COL[8953] = 1'b0;
assign COL[8954] = 1'b0;
assign COL[8955] = 1'b0;
assign COL[8956] = 1'b0;
assign COL[8957] = 1'b0;
assign COL[8958] = 1'b0;
assign COL[8959] = 1'b0;
assign COL[8960] = 1'b0;
assign COL[8961] = 1'b1;
assign COL[8962] = 1'b1;
assign COL[8963] = 1'b1;
assign COL[8964] = 1'b1;
assign COL[8965] = 1'b1;
assign COL[8966] = 1'b0;
assign COL[8967] = 1'b0;
assign COL[8968] = 1'b0;
assign COL[8969] = 1'b0;
assign COL[8970] = 1'b0;
assign COL[8971] = 1'b0;
assign COL[8972] = 1'b0;
assign COL[8973] = 1'b0;
assign COL[8974] = 1'b0;
assign COL[8975] = 1'b0;
assign COL[8976] = 1'b0;
assign COL[8977] = 1'b0;
assign COL[8978] = 1'b0;
assign COL[8979] = 1'b0;
assign COL[8980] = 1'b0;
assign COL[8981] = 1'b0;
assign COL[8982] = 1'b0;
assign COL[8983] = 1'b0;
assign COL[8984] = 1'b0;
assign COL[8985] = 1'b0;
assign COL[8986] = 1'b0;
assign COL[8987] = 1'b0;
assign COL[8988] = 1'b0;
assign COL[8989] = 1'b1;
assign COL[8990] = 1'b1;
assign COL[8991] = 1'b1;
assign COL[8992] = 1'b1;
assign COL[8993] = 1'b0;
assign COL[8994] = 1'b0;
assign COL[8995] = 1'b0;
assign COL[8996] = 1'b0;
assign COL[8997] = 1'b0;
assign COL[8998] = 1'b0;
assign COL[8999] = 1'b0;
assign COL[9000] = 1'b0;
assign COL[9001] = 1'b0;
assign COL[9002] = 1'b0;
assign COL[9003] = 1'b0;
assign COL[9004] = 1'b0;
assign COL[9005] = 1'b0;
assign COL[9006] = 1'b0;
assign COL[9007] = 1'b0;
assign COL[9008] = 1'b0;
assign COL[9009] = 1'b0;
assign COL[9010] = 1'b0;
assign COL[9011] = 1'b0;
assign COL[9012] = 1'b0;
assign COL[9013] = 1'b0;
assign COL[9014] = 1'b0;
assign COL[9015] = 1'b0;
assign COL[9016] = 1'b0;
assign COL[9017] = 1'b0;
assign COL[9018] = 1'b1;
assign COL[9019] = 1'b1;
assign COL[9020] = 1'b1;
assign COL[9021] = 1'b1;
assign COL[9022] = 1'b0;
assign COL[9023] = 1'b0;
assign COL[9024] = 1'b0;
assign COL[9025] = 1'b0;
assign COL[9026] = 1'b0;
assign COL[9027] = 1'b0;
assign COL[9028] = 1'b0;
assign COL[9029] = 1'b0;
assign COL[9030] = 1'b1;
assign COL[9031] = 1'b1;
assign COL[9032] = 1'b1;
assign COL[9033] = 1'b1;
assign COL[9034] = 1'b1;
assign COL[9035] = 1'b0;
assign COL[9036] = 1'b0;
assign COL[9037] = 1'b0;
assign COL[9038] = 1'b0;
assign COL[9039] = 1'b0;
assign COL[9040] = 1'b0;
assign COL[9041] = 1'b0;
assign COL[9042] = 1'b0;
assign COL[9043] = 1'b0;
assign COL[9044] = 1'b0;
assign COL[9045] = 1'b0;
assign COL[9046] = 1'b0;
assign COL[9047] = 1'b0;
assign COL[9048] = 1'b0;
assign COL[9049] = 1'b0;
assign COL[9050] = 1'b1;
assign COL[9051] = 1'b1;
assign COL[9052] = 1'b1;
assign COL[9053] = 1'b1;
assign COL[9054] = 1'b1;
assign COL[9055] = 1'b0;
assign COL[9056] = 1'b0;
assign COL[9057] = 1'b0;
assign COL[9058] = 1'b0;
assign COL[9059] = 1'b0;
assign COL[9060] = 1'b0;
assign COL[9061] = 1'b0;
assign COL[9062] = 1'b0;
assign COL[9063] = 1'b0;
assign COL[9064] = 1'b0;
assign COL[9065] = 1'b0;
assign COL[9066] = 1'b0;
assign COL[9067] = 1'b0;
assign COL[9068] = 1'b0;
assign COL[9069] = 1'b0;
assign COL[9070] = 1'b0;
assign COL[9071] = 1'b0;
assign COL[9072] = 1'b0;
assign COL[9073] = 1'b0;
assign COL[9074] = 1'b0;
assign COL[9075] = 1'b0;
assign COL[9076] = 1'b0;
assign COL[9077] = 1'b0;
assign COL[9078] = 1'b0;
assign COL[9079] = 1'b0;
assign COL[9080] = 1'b0;
assign COL[9081] = 1'b0;
assign COL[9082] = 1'b0;
assign COL[9083] = 1'b0;
assign COL[9084] = 1'b0;
assign COL[9085] = 1'b0;
assign COL[9086] = 1'b0;
assign COL[9087] = 1'b0;
assign COL[9088] = 1'b0;
assign COL[9089] = 1'b0;
assign COL[9090] = 1'b0;
assign COL[9091] = 1'b0;
assign COL[9092] = 1'b0;
assign COL[9093] = 1'b0;
assign COL[9094] = 1'b0;
assign COL[9095] = 1'b0;
assign COL[9096] = 1'b0;
assign COL[9097] = 1'b0;
assign COL[9098] = 1'b0;
assign COL[9099] = 1'b0;
assign COL[9100] = 1'b0;
assign COL[9101] = 1'b0;
assign COL[9102] = 1'b0;
assign COL[9103] = 1'b0;
assign COL[9104] = 1'b0;
assign COL[9105] = 1'b0;
assign COL[9106] = 1'b0;
assign COL[9107] = 1'b0;
assign COL[9108] = 1'b0;
assign COL[9109] = 1'b0;
assign COL[9110] = 1'b0;
assign COL[9111] = 1'b0;
assign COL[9112] = 1'b0;
assign COL[9113] = 1'b0;
assign COL[9114] = 1'b0;
assign COL[9115] = 1'b0;
assign COL[9116] = 1'b0;
assign COL[9117] = 1'b0;
assign COL[9118] = 1'b0;
assign COL[9119] = 1'b0;
assign COL[9120] = 1'b0;
assign COL[9121] = 1'b1;
assign COL[9122] = 1'b1;
assign COL[9123] = 1'b1;
assign COL[9124] = 1'b1;
assign COL[9125] = 1'b1;
assign COL[9126] = 1'b0;
assign COL[9127] = 1'b0;
assign COL[9128] = 1'b0;
assign COL[9129] = 1'b0;
assign COL[9130] = 1'b0;
assign COL[9131] = 1'b0;
assign COL[9132] = 1'b0;
assign COL[9133] = 1'b0;
assign COL[9134] = 1'b0;
assign COL[9135] = 1'b0;
assign COL[9136] = 1'b0;
assign COL[9137] = 1'b0;
assign COL[9138] = 1'b0;
assign COL[9139] = 1'b0;
assign COL[9140] = 1'b0;
assign COL[9141] = 1'b0;
assign COL[9142] = 1'b0;
assign COL[9143] = 1'b0;
assign COL[9144] = 1'b0;
assign COL[9145] = 1'b0;
assign COL[9146] = 1'b0;
assign COL[9147] = 1'b0;
assign COL[9148] = 1'b0;
assign COL[9149] = 1'b1;
assign COL[9150] = 1'b1;
assign COL[9151] = 1'b1;
assign COL[9152] = 1'b1;
assign COL[9153] = 1'b0;
assign COL[9154] = 1'b0;
assign COL[9155] = 1'b0;
assign COL[9156] = 1'b0;
assign COL[9157] = 1'b0;
assign COL[9158] = 1'b0;
assign COL[9159] = 1'b0;
assign COL[9160] = 1'b0;
assign COL[9161] = 1'b0;
assign COL[9162] = 1'b0;
assign COL[9163] = 1'b0;
assign COL[9164] = 1'b0;
assign COL[9165] = 1'b0;
assign COL[9166] = 1'b0;
assign COL[9167] = 1'b0;
assign COL[9168] = 1'b0;
assign COL[9169] = 1'b0;
assign COL[9170] = 1'b0;
assign COL[9171] = 1'b0;
assign COL[9172] = 1'b0;
assign COL[9173] = 1'b0;
assign COL[9174] = 1'b0;
assign COL[9175] = 1'b0;
assign COL[9176] = 1'b0;
assign COL[9177] = 1'b0;
assign COL[9178] = 1'b1;
assign COL[9179] = 1'b1;
assign COL[9180] = 1'b1;
assign COL[9181] = 1'b1;
assign COL[9182] = 1'b0;
assign COL[9183] = 1'b0;
assign COL[9184] = 1'b0;
assign COL[9185] = 1'b0;
assign COL[9186] = 1'b0;
assign COL[9187] = 1'b0;
assign COL[9188] = 1'b0;
assign COL[9189] = 1'b0;
assign COL[9190] = 1'b1;
assign COL[9191] = 1'b1;
assign COL[9192] = 1'b1;
assign COL[9193] = 1'b1;
assign COL[9194] = 1'b1;
assign COL[9195] = 1'b0;
assign COL[9196] = 1'b0;
assign COL[9197] = 1'b0;
assign COL[9198] = 1'b0;
assign COL[9199] = 1'b0;
assign COL[9200] = 1'b0;
assign COL[9201] = 1'b0;
assign COL[9202] = 1'b0;
assign COL[9203] = 1'b0;
assign COL[9204] = 1'b0;
assign COL[9205] = 1'b0;
assign COL[9206] = 1'b0;
assign COL[9207] = 1'b0;
assign COL[9208] = 1'b0;
assign COL[9209] = 1'b0;
assign COL[9210] = 1'b1;
assign COL[9211] = 1'b1;
assign COL[9212] = 1'b1;
assign COL[9213] = 1'b1;
assign COL[9214] = 1'b1;
assign COL[9215] = 1'b0;
assign COL[9216] = 1'b0;
assign COL[9217] = 1'b0;
assign COL[9218] = 1'b0;
assign COL[9219] = 1'b0;
assign COL[9220] = 1'b0;
assign COL[9221] = 1'b0;
assign COL[9222] = 1'b0;
assign COL[9223] = 1'b0;
assign COL[9224] = 1'b0;
assign COL[9225] = 1'b0;
assign COL[9226] = 1'b0;
assign COL[9227] = 1'b0;
assign COL[9228] = 1'b0;
assign COL[9229] = 1'b0;
assign COL[9230] = 1'b0;
assign COL[9231] = 1'b0;
assign COL[9232] = 1'b0;
assign COL[9233] = 1'b0;
assign COL[9234] = 1'b0;
assign COL[9235] = 1'b0;
assign COL[9236] = 1'b0;
assign COL[9237] = 1'b0;
assign COL[9238] = 1'b0;
assign COL[9239] = 1'b0;
assign COL[9240] = 1'b0;
assign COL[9241] = 1'b0;
assign COL[9242] = 1'b0;
assign COL[9243] = 1'b0;
assign COL[9244] = 1'b0;
assign COL[9245] = 1'b0;
assign COL[9246] = 1'b0;
assign COL[9247] = 1'b0;
assign COL[9248] = 1'b0;
assign COL[9249] = 1'b0;
assign COL[9250] = 1'b0;
assign COL[9251] = 1'b0;
assign COL[9252] = 1'b0;
assign COL[9253] = 1'b0;
assign COL[9254] = 1'b0;
assign COL[9255] = 1'b0;
assign COL[9256] = 1'b0;
assign COL[9257] = 1'b0;
assign COL[9258] = 1'b0;
assign COL[9259] = 1'b0;
assign COL[9260] = 1'b0;
assign COL[9261] = 1'b0;
assign COL[9262] = 1'b0;
assign COL[9263] = 1'b0;
assign COL[9264] = 1'b0;
assign COL[9265] = 1'b0;
assign COL[9266] = 1'b0;
assign COL[9267] = 1'b0;
assign COL[9268] = 1'b0;
assign COL[9269] = 1'b0;
assign COL[9270] = 1'b0;
assign COL[9271] = 1'b0;
assign COL[9272] = 1'b0;
assign COL[9273] = 1'b0;
assign COL[9274] = 1'b0;
assign COL[9275] = 1'b0;
assign COL[9276] = 1'b0;
assign COL[9277] = 1'b0;
assign COL[9278] = 1'b0;
assign COL[9279] = 1'b0;
assign COL[9280] = 1'b0;
assign COL[9281] = 1'b1;
assign COL[9282] = 1'b1;
assign COL[9283] = 1'b1;
assign COL[9284] = 1'b1;
assign COL[9285] = 1'b1;
assign COL[9286] = 1'b0;
assign COL[9287] = 1'b0;
assign COL[9288] = 1'b0;
assign COL[9289] = 1'b0;
assign COL[9290] = 1'b0;
assign COL[9291] = 1'b0;
assign COL[9292] = 1'b0;
assign COL[9293] = 1'b0;
assign COL[9294] = 1'b0;
assign COL[9295] = 1'b0;
assign COL[9296] = 1'b0;
assign COL[9297] = 1'b0;
assign COL[9298] = 1'b0;
assign COL[9299] = 1'b0;
assign COL[9300] = 1'b0;
assign COL[9301] = 1'b0;
assign COL[9302] = 1'b0;
assign COL[9303] = 1'b0;
assign COL[9304] = 1'b0;
assign COL[9305] = 1'b0;
assign COL[9306] = 1'b0;
assign COL[9307] = 1'b0;
assign COL[9308] = 1'b0;
assign COL[9309] = 1'b1;
assign COL[9310] = 1'b1;
assign COL[9311] = 1'b1;
assign COL[9312] = 1'b1;
assign COL[9313] = 1'b0;
assign COL[9314] = 1'b0;
assign COL[9315] = 1'b0;
assign COL[9316] = 1'b0;
assign COL[9317] = 1'b0;
assign COL[9318] = 1'b0;
assign COL[9319] = 1'b0;
assign COL[9320] = 1'b0;
assign COL[9321] = 1'b0;
assign COL[9322] = 1'b0;
assign COL[9323] = 1'b0;
assign COL[9324] = 1'b0;
assign COL[9325] = 1'b0;
assign COL[9326] = 1'b0;
assign COL[9327] = 1'b0;
assign COL[9328] = 1'b0;
assign COL[9329] = 1'b0;
assign COL[9330] = 1'b0;
assign COL[9331] = 1'b0;
assign COL[9332] = 1'b0;
assign COL[9333] = 1'b0;
assign COL[9334] = 1'b0;
assign COL[9335] = 1'b0;
assign COL[9336] = 1'b0;
assign COL[9337] = 1'b0;
assign COL[9338] = 1'b1;
assign COL[9339] = 1'b1;
assign COL[9340] = 1'b1;
assign COL[9341] = 1'b1;
assign COL[9342] = 1'b0;
assign COL[9343] = 1'b0;
assign COL[9344] = 1'b0;
assign COL[9345] = 1'b0;
assign COL[9346] = 1'b0;
assign COL[9347] = 1'b0;
assign COL[9348] = 1'b0;
assign COL[9349] = 1'b0;
assign COL[9350] = 1'b1;
assign COL[9351] = 1'b1;
assign COL[9352] = 1'b1;
assign COL[9353] = 1'b1;
assign COL[9354] = 1'b1;
assign COL[9355] = 1'b0;
assign COL[9356] = 1'b0;
assign COL[9357] = 1'b0;
assign COL[9358] = 1'b0;
assign COL[9359] = 1'b0;
assign COL[9360] = 1'b0;
assign COL[9361] = 1'b0;
assign COL[9362] = 1'b0;
assign COL[9363] = 1'b0;
assign COL[9364] = 1'b0;
assign COL[9365] = 1'b0;
assign COL[9366] = 1'b0;
assign COL[9367] = 1'b0;
assign COL[9368] = 1'b0;
assign COL[9369] = 1'b0;
assign COL[9370] = 1'b1;
assign COL[9371] = 1'b1;
assign COL[9372] = 1'b1;
assign COL[9373] = 1'b1;
assign COL[9374] = 1'b1;
assign COL[9375] = 1'b0;
assign COL[9376] = 1'b0;
assign COL[9377] = 1'b0;
assign COL[9378] = 1'b0;
assign COL[9379] = 1'b0;
assign COL[9380] = 1'b0;
assign COL[9381] = 1'b0;
assign COL[9382] = 1'b0;
assign COL[9383] = 1'b0;
assign COL[9384] = 1'b0;
assign COL[9385] = 1'b0;
assign COL[9386] = 1'b0;
assign COL[9387] = 1'b0;
assign COL[9388] = 1'b0;
assign COL[9389] = 1'b0;
assign COL[9390] = 1'b0;
assign COL[9391] = 1'b0;
assign COL[9392] = 1'b0;
assign COL[9393] = 1'b0;
assign COL[9394] = 1'b0;
assign COL[9395] = 1'b0;
assign COL[9396] = 1'b0;
assign COL[9397] = 1'b0;
assign COL[9398] = 1'b0;
assign COL[9399] = 1'b0;
assign COL[9400] = 1'b0;
assign COL[9401] = 1'b0;
assign COL[9402] = 1'b0;
assign COL[9403] = 1'b0;
assign COL[9404] = 1'b0;
assign COL[9405] = 1'b0;
assign COL[9406] = 1'b0;
assign COL[9407] = 1'b0;
assign COL[9408] = 1'b0;
assign COL[9409] = 1'b0;
assign COL[9410] = 1'b0;
assign COL[9411] = 1'b0;
assign COL[9412] = 1'b0;
assign COL[9413] = 1'b0;
assign COL[9414] = 1'b0;
assign COL[9415] = 1'b0;
assign COL[9416] = 1'b0;
assign COL[9417] = 1'b0;
assign COL[9418] = 1'b0;
assign COL[9419] = 1'b0;
assign COL[9420] = 1'b0;
assign COL[9421] = 1'b0;
assign COL[9422] = 1'b0;
assign COL[9423] = 1'b0;
assign COL[9424] = 1'b0;
assign COL[9425] = 1'b0;
assign COL[9426] = 1'b0;
assign COL[9427] = 1'b0;
assign COL[9428] = 1'b0;
assign COL[9429] = 1'b0;
assign COL[9430] = 1'b0;
assign COL[9431] = 1'b0;
assign COL[9432] = 1'b0;
assign COL[9433] = 1'b0;
assign COL[9434] = 1'b0;
assign COL[9435] = 1'b0;
assign COL[9436] = 1'b0;
assign COL[9437] = 1'b0;
assign COL[9438] = 1'b0;
assign COL[9439] = 1'b0;
assign COL[9440] = 1'b0;
assign COL[9441] = 1'b1;
assign COL[9442] = 1'b1;
assign COL[9443] = 1'b1;
assign COL[9444] = 1'b1;
assign COL[9445] = 1'b1;
assign COL[9446] = 1'b0;
assign COL[9447] = 1'b0;
assign COL[9448] = 1'b0;
assign COL[9449] = 1'b0;
assign COL[9450] = 1'b0;
assign COL[9451] = 1'b0;
assign COL[9452] = 1'b0;
assign COL[9453] = 1'b0;
assign COL[9454] = 1'b0;
assign COL[9455] = 1'b0;
assign COL[9456] = 1'b0;
assign COL[9457] = 1'b0;
assign COL[9458] = 1'b0;
assign COL[9459] = 1'b0;
assign COL[9460] = 1'b0;
assign COL[9461] = 1'b0;
assign COL[9462] = 1'b0;
assign COL[9463] = 1'b0;
assign COL[9464] = 1'b0;
assign COL[9465] = 1'b0;
assign COL[9466] = 1'b0;
assign COL[9467] = 1'b0;
assign COL[9468] = 1'b0;
assign COL[9469] = 1'b1;
assign COL[9470] = 1'b1;
assign COL[9471] = 1'b1;
assign COL[9472] = 1'b1;
assign COL[9473] = 1'b0;
assign COL[9474] = 1'b0;
assign COL[9475] = 1'b0;
assign COL[9476] = 1'b0;
assign COL[9477] = 1'b0;
assign COL[9478] = 1'b0;
assign COL[9479] = 1'b0;
assign COL[9480] = 1'b0;
assign COL[9481] = 1'b0;
assign COL[9482] = 1'b0;
assign COL[9483] = 1'b0;
assign COL[9484] = 1'b0;
assign COL[9485] = 1'b0;
assign COL[9486] = 1'b0;
assign COL[9487] = 1'b0;
assign COL[9488] = 1'b0;
assign COL[9489] = 1'b0;
assign COL[9490] = 1'b0;
assign COL[9491] = 1'b0;
assign COL[9492] = 1'b0;
assign COL[9493] = 1'b0;
assign COL[9494] = 1'b0;
assign COL[9495] = 1'b0;
assign COL[9496] = 1'b0;
assign COL[9497] = 1'b0;
assign COL[9498] = 1'b1;
assign COL[9499] = 1'b1;
assign COL[9500] = 1'b1;
assign COL[9501] = 1'b1;
assign COL[9502] = 1'b0;
assign COL[9503] = 1'b0;
assign COL[9504] = 1'b0;
assign COL[9505] = 1'b0;
assign COL[9506] = 1'b0;
assign COL[9507] = 1'b0;
assign COL[9508] = 1'b0;
assign COL[9509] = 1'b0;
assign COL[9510] = 1'b1;
assign COL[9511] = 1'b1;
assign COL[9512] = 1'b1;
assign COL[9513] = 1'b1;
assign COL[9514] = 1'b1;
assign COL[9515] = 1'b0;
assign COL[9516] = 1'b0;
assign COL[9517] = 1'b0;
assign COL[9518] = 1'b0;
assign COL[9519] = 1'b0;
assign COL[9520] = 1'b0;
assign COL[9521] = 1'b0;
assign COL[9522] = 1'b0;
assign COL[9523] = 1'b0;
assign COL[9524] = 1'b0;
assign COL[9525] = 1'b0;
assign COL[9526] = 1'b0;
assign COL[9527] = 1'b0;
assign COL[9528] = 1'b0;
assign COL[9529] = 1'b0;
assign COL[9530] = 1'b1;
assign COL[9531] = 1'b1;
assign COL[9532] = 1'b1;
assign COL[9533] = 1'b1;
assign COL[9534] = 1'b1;
assign COL[9535] = 1'b0;
assign COL[9536] = 1'b0;
assign COL[9537] = 1'b0;
assign COL[9538] = 1'b0;
assign COL[9539] = 1'b0;
assign COL[9540] = 1'b0;
assign COL[9541] = 1'b0;
assign COL[9542] = 1'b0;
assign COL[9543] = 1'b0;
assign COL[9544] = 1'b0;
assign COL[9545] = 1'b0;
assign COL[9546] = 1'b0;
assign COL[9547] = 1'b0;
assign COL[9548] = 1'b0;
assign COL[9549] = 1'b0;
assign COL[9550] = 1'b0;
assign COL[9551] = 1'b0;
assign COL[9552] = 1'b0;
assign COL[9553] = 1'b0;
assign COL[9554] = 1'b0;
assign COL[9555] = 1'b0;
assign COL[9556] = 1'b0;
assign COL[9557] = 1'b0;
assign COL[9558] = 1'b0;
assign COL[9559] = 1'b0;
assign COL[9560] = 1'b0;
assign COL[9561] = 1'b0;
assign COL[9562] = 1'b0;
assign COL[9563] = 1'b0;
assign COL[9564] = 1'b0;
assign COL[9565] = 1'b0;
assign COL[9566] = 1'b0;
assign COL[9567] = 1'b0;
assign COL[9568] = 1'b0;
assign COL[9569] = 1'b0;
assign COL[9570] = 1'b0;
assign COL[9571] = 1'b0;
assign COL[9572] = 1'b0;
assign COL[9573] = 1'b0;
assign COL[9574] = 1'b0;
assign COL[9575] = 1'b0;
assign COL[9576] = 1'b0;
assign COL[9577] = 1'b0;
assign COL[9578] = 1'b0;
assign COL[9579] = 1'b0;
assign COL[9580] = 1'b0;
assign COL[9581] = 1'b0;
assign COL[9582] = 1'b0;
assign COL[9583] = 1'b0;
assign COL[9584] = 1'b0;
assign COL[9585] = 1'b0;
assign COL[9586] = 1'b0;
assign COL[9587] = 1'b0;
assign COL[9588] = 1'b0;
assign COL[9589] = 1'b0;
assign COL[9590] = 1'b0;
assign COL[9591] = 1'b0;
assign COL[9592] = 1'b0;
assign COL[9593] = 1'b0;
assign COL[9594] = 1'b0;
assign COL[9595] = 1'b0;
assign COL[9596] = 1'b0;
assign COL[9597] = 1'b0;
assign COL[9598] = 1'b0;
assign COL[9599] = 1'b0;
assign COL[9600] = 1'b0;
assign COL[9601] = 1'b1;
assign COL[9602] = 1'b1;
assign COL[9603] = 1'b1;
assign COL[9604] = 1'b1;
assign COL[9605] = 1'b1;
assign COL[9606] = 1'b0;
assign COL[9607] = 1'b0;
assign COL[9608] = 1'b0;
assign COL[9609] = 1'b0;
assign COL[9610] = 1'b0;
assign COL[9611] = 1'b0;
assign COL[9612] = 1'b0;
assign COL[9613] = 1'b0;
assign COL[9614] = 1'b0;
assign COL[9615] = 1'b0;
assign COL[9616] = 1'b0;
assign COL[9617] = 1'b0;
assign COL[9618] = 1'b0;
assign COL[9619] = 1'b0;
assign COL[9620] = 1'b0;
assign COL[9621] = 1'b0;
assign COL[9622] = 1'b0;
assign COL[9623] = 1'b0;
assign COL[9624] = 1'b0;
assign COL[9625] = 1'b0;
assign COL[9626] = 1'b0;
assign COL[9627] = 1'b0;
assign COL[9628] = 1'b0;
assign COL[9629] = 1'b1;
assign COL[9630] = 1'b1;
assign COL[9631] = 1'b1;
assign COL[9632] = 1'b1;
assign COL[9633] = 1'b0;
assign COL[9634] = 1'b0;
assign COL[9635] = 1'b0;
assign COL[9636] = 1'b0;
assign COL[9637] = 1'b0;
assign COL[9638] = 1'b0;
assign COL[9639] = 1'b0;
assign COL[9640] = 1'b0;
assign COL[9641] = 1'b0;
assign COL[9642] = 1'b0;
assign COL[9643] = 1'b0;
assign COL[9644] = 1'b0;
assign COL[9645] = 1'b0;
assign COL[9646] = 1'b0;
assign COL[9647] = 1'b0;
assign COL[9648] = 1'b0;
assign COL[9649] = 1'b0;
assign COL[9650] = 1'b0;
assign COL[9651] = 1'b0;
assign COL[9652] = 1'b0;
assign COL[9653] = 1'b0;
assign COL[9654] = 1'b0;
assign COL[9655] = 1'b0;
assign COL[9656] = 1'b0;
assign COL[9657] = 1'b0;
assign COL[9658] = 1'b1;
assign COL[9659] = 1'b1;
assign COL[9660] = 1'b1;
assign COL[9661] = 1'b1;
assign COL[9662] = 1'b0;
assign COL[9663] = 1'b0;
assign COL[9664] = 1'b0;
assign COL[9665] = 1'b0;
assign COL[9666] = 1'b0;
assign COL[9667] = 1'b0;
assign COL[9668] = 1'b0;
assign COL[9669] = 1'b0;
assign COL[9670] = 1'b1;
assign COL[9671] = 1'b1;
assign COL[9672] = 1'b1;
assign COL[9673] = 1'b1;
assign COL[9674] = 1'b1;
assign COL[9675] = 1'b0;
assign COL[9676] = 1'b0;
assign COL[9677] = 1'b0;
assign COL[9678] = 1'b0;
assign COL[9679] = 1'b0;
assign COL[9680] = 1'b0;
assign COL[9681] = 1'b0;
assign COL[9682] = 1'b0;
assign COL[9683] = 1'b0;
assign COL[9684] = 1'b0;
assign COL[9685] = 1'b0;
assign COL[9686] = 1'b0;
assign COL[9687] = 1'b0;
assign COL[9688] = 1'b0;
assign COL[9689] = 1'b0;
assign COL[9690] = 1'b1;
assign COL[9691] = 1'b1;
assign COL[9692] = 1'b1;
assign COL[9693] = 1'b1;
assign COL[9694] = 1'b1;
assign COL[9695] = 1'b0;
assign COL[9696] = 1'b0;
assign COL[9697] = 1'b0;
assign COL[9698] = 1'b0;
assign COL[9699] = 1'b0;
assign COL[9700] = 1'b0;
assign COL[9701] = 1'b0;
assign COL[9702] = 1'b0;
assign COL[9703] = 1'b0;
assign COL[9704] = 1'b0;
assign COL[9705] = 1'b0;
assign COL[9706] = 1'b0;
assign COL[9707] = 1'b0;
assign COL[9708] = 1'b0;
assign COL[9709] = 1'b0;
assign COL[9710] = 1'b0;
assign COL[9711] = 1'b0;
assign COL[9712] = 1'b0;
assign COL[9713] = 1'b0;
assign COL[9714] = 1'b0;
assign COL[9715] = 1'b0;
assign COL[9716] = 1'b0;
assign COL[9717] = 1'b0;
assign COL[9718] = 1'b0;
assign COL[9719] = 1'b0;
assign COL[9720] = 1'b0;
assign COL[9721] = 1'b0;
assign COL[9722] = 1'b0;
assign COL[9723] = 1'b0;
assign COL[9724] = 1'b0;
assign COL[9725] = 1'b0;
assign COL[9726] = 1'b0;
assign COL[9727] = 1'b0;
assign COL[9728] = 1'b0;
assign COL[9729] = 1'b0;
assign COL[9730] = 1'b0;
assign COL[9731] = 1'b0;
assign COL[9732] = 1'b0;
assign COL[9733] = 1'b0;
assign COL[9734] = 1'b0;
assign COL[9735] = 1'b0;
assign COL[9736] = 1'b0;
assign COL[9737] = 1'b0;
assign COL[9738] = 1'b0;
assign COL[9739] = 1'b0;
assign COL[9740] = 1'b0;
assign COL[9741] = 1'b0;
assign COL[9742] = 1'b0;
assign COL[9743] = 1'b0;
assign COL[9744] = 1'b0;
assign COL[9745] = 1'b0;
assign COL[9746] = 1'b0;
assign COL[9747] = 1'b0;
assign COL[9748] = 1'b0;
assign COL[9749] = 1'b0;
assign COL[9750] = 1'b0;
assign COL[9751] = 1'b0;
assign COL[9752] = 1'b0;
assign COL[9753] = 1'b0;
assign COL[9754] = 1'b0;
assign COL[9755] = 1'b0;
assign COL[9756] = 1'b0;
assign COL[9757] = 1'b0;
assign COL[9758] = 1'b0;
assign COL[9759] = 1'b0;
assign COL[9760] = 1'b0;
assign COL[9761] = 1'b1;
assign COL[9762] = 1'b1;
assign COL[9763] = 1'b1;
assign COL[9764] = 1'b1;
assign COL[9765] = 1'b1;
assign COL[9766] = 1'b0;
assign COL[9767] = 1'b0;
assign COL[9768] = 1'b0;
assign COL[9769] = 1'b0;
assign COL[9770] = 1'b0;
assign COL[9771] = 1'b0;
assign COL[9772] = 1'b0;
assign COL[9773] = 1'b0;
assign COL[9774] = 1'b0;
assign COL[9775] = 1'b0;
assign COL[9776] = 1'b0;
assign COL[9777] = 1'b0;
assign COL[9778] = 1'b0;
assign COL[9779] = 1'b0;
assign COL[9780] = 1'b0;
assign COL[9781] = 1'b0;
assign COL[9782] = 1'b0;
assign COL[9783] = 1'b0;
assign COL[9784] = 1'b0;
assign COL[9785] = 1'b0;
assign COL[9786] = 1'b0;
assign COL[9787] = 1'b0;
assign COL[9788] = 1'b0;
assign COL[9789] = 1'b1;
assign COL[9790] = 1'b1;
assign COL[9791] = 1'b1;
assign COL[9792] = 1'b1;
assign COL[9793] = 1'b0;
assign COL[9794] = 1'b0;
assign COL[9795] = 1'b0;
assign COL[9796] = 1'b0;
assign COL[9797] = 1'b0;
assign COL[9798] = 1'b0;
assign COL[9799] = 1'b0;
assign COL[9800] = 1'b0;
assign COL[9801] = 1'b0;
assign COL[9802] = 1'b0;
assign COL[9803] = 1'b0;
assign COL[9804] = 1'b0;
assign COL[9805] = 1'b0;
assign COL[9806] = 1'b0;
assign COL[9807] = 1'b0;
assign COL[9808] = 1'b0;
assign COL[9809] = 1'b0;
assign COL[9810] = 1'b0;
assign COL[9811] = 1'b0;
assign COL[9812] = 1'b0;
assign COL[9813] = 1'b0;
assign COL[9814] = 1'b0;
assign COL[9815] = 1'b0;
assign COL[9816] = 1'b0;
assign COL[9817] = 1'b0;
assign COL[9818] = 1'b1;
assign COL[9819] = 1'b1;
assign COL[9820] = 1'b1;
assign COL[9821] = 1'b1;
assign COL[9822] = 1'b0;
assign COL[9823] = 1'b0;
assign COL[9824] = 1'b0;
assign COL[9825] = 1'b0;
assign COL[9826] = 1'b0;
assign COL[9827] = 1'b0;
assign COL[9828] = 1'b0;
assign COL[9829] = 1'b0;
assign COL[9830] = 1'b1;
assign COL[9831] = 1'b1;
assign COL[9832] = 1'b1;
assign COL[9833] = 1'b1;
assign COL[9834] = 1'b1;
assign COL[9835] = 1'b1;
assign COL[9836] = 1'b1;
assign COL[9837] = 1'b1;
assign COL[9838] = 1'b1;
assign COL[9839] = 1'b1;
assign COL[9840] = 1'b1;
assign COL[9841] = 1'b1;
assign COL[9842] = 1'b1;
assign COL[9843] = 1'b1;
assign COL[9844] = 1'b1;
assign COL[9845] = 1'b1;
assign COL[9846] = 1'b1;
assign COL[9847] = 1'b1;
assign COL[9848] = 1'b1;
assign COL[9849] = 1'b1;
assign COL[9850] = 1'b1;
assign COL[9851] = 1'b1;
assign COL[9852] = 1'b1;
assign COL[9853] = 1'b1;
assign COL[9854] = 1'b1;
assign COL[9855] = 1'b0;
assign COL[9856] = 1'b0;
assign COL[9857] = 1'b0;
assign COL[9858] = 1'b0;
assign COL[9859] = 1'b0;
assign COL[9860] = 1'b0;
assign COL[9861] = 1'b0;
assign COL[9862] = 1'b0;
assign COL[9863] = 1'b0;
assign COL[9864] = 1'b0;
assign COL[9865] = 1'b0;
assign COL[9866] = 1'b0;
assign COL[9867] = 1'b0;
assign COL[9868] = 1'b0;
assign COL[9869] = 1'b0;
assign COL[9870] = 1'b0;
assign COL[9871] = 1'b0;
assign COL[9872] = 1'b0;
assign COL[9873] = 1'b0;
assign COL[9874] = 1'b0;
assign COL[9875] = 1'b0;
assign COL[9876] = 1'b0;
assign COL[9877] = 1'b0;
assign COL[9878] = 1'b0;
assign COL[9879] = 1'b0;
assign COL[9880] = 1'b0;
assign COL[9881] = 1'b0;
assign COL[9882] = 1'b0;
assign COL[9883] = 1'b0;
assign COL[9884] = 1'b0;
assign COL[9885] = 1'b0;
assign COL[9886] = 1'b0;
assign COL[9887] = 1'b0;
assign COL[9888] = 1'b0;
assign COL[9889] = 1'b0;
assign COL[9890] = 1'b0;
assign COL[9891] = 1'b0;
assign COL[9892] = 1'b0;
assign COL[9893] = 1'b0;
assign COL[9894] = 1'b0;
assign COL[9895] = 1'b0;
assign COL[9896] = 1'b0;
assign COL[9897] = 1'b0;
assign COL[9898] = 1'b0;
assign COL[9899] = 1'b0;
assign COL[9900] = 1'b0;
assign COL[9901] = 1'b0;
assign COL[9902] = 1'b0;
assign COL[9903] = 1'b0;
assign COL[9904] = 1'b0;
assign COL[9905] = 1'b0;
assign COL[9906] = 1'b0;
assign COL[9907] = 1'b0;
assign COL[9908] = 1'b0;
assign COL[9909] = 1'b0;
assign COL[9910] = 1'b0;
assign COL[9911] = 1'b0;
assign COL[9912] = 1'b0;
assign COL[9913] = 1'b0;
assign COL[9914] = 1'b0;
assign COL[9915] = 1'b0;
assign COL[9916] = 1'b0;
assign COL[9917] = 1'b0;
assign COL[9918] = 1'b0;
assign COL[9919] = 1'b0;
assign COL[9920] = 1'b0;
assign COL[9921] = 1'b1;
assign COL[9922] = 1'b1;
assign COL[9923] = 1'b1;
assign COL[9924] = 1'b1;
assign COL[9925] = 1'b1;
assign COL[9926] = 1'b0;
assign COL[9927] = 1'b0;
assign COL[9928] = 1'b0;
assign COL[9929] = 1'b0;
assign COL[9930] = 1'b0;
assign COL[9931] = 1'b0;
assign COL[9932] = 1'b0;
assign COL[9933] = 1'b0;
assign COL[9934] = 1'b0;
assign COL[9935] = 1'b0;
assign COL[9936] = 1'b0;
assign COL[9937] = 1'b0;
assign COL[9938] = 1'b0;
assign COL[9939] = 1'b0;
assign COL[9940] = 1'b0;
assign COL[9941] = 1'b0;
assign COL[9942] = 1'b0;
assign COL[9943] = 1'b0;
assign COL[9944] = 1'b0;
assign COL[9945] = 1'b0;
assign COL[9946] = 1'b0;
assign COL[9947] = 1'b0;
assign COL[9948] = 1'b0;
assign COL[9949] = 1'b1;
assign COL[9950] = 1'b1;
assign COL[9951] = 1'b1;
assign COL[9952] = 1'b1;
assign COL[9953] = 1'b0;
assign COL[9954] = 1'b0;
assign COL[9955] = 1'b0;
assign COL[9956] = 1'b0;
assign COL[9957] = 1'b0;
assign COL[9958] = 1'b0;
assign COL[9959] = 1'b0;
assign COL[9960] = 1'b0;
assign COL[9961] = 1'b0;
assign COL[9962] = 1'b0;
assign COL[9963] = 1'b0;
assign COL[9964] = 1'b0;
assign COL[9965] = 1'b1;
assign COL[9966] = 1'b1;
assign COL[9967] = 1'b1;
assign COL[9968] = 1'b1;
assign COL[9969] = 1'b1;
assign COL[9970] = 1'b1;
assign COL[9971] = 1'b1;
assign COL[9972] = 1'b1;
assign COL[9973] = 1'b1;
assign COL[9974] = 1'b1;
assign COL[9975] = 1'b1;
assign COL[9976] = 1'b1;
assign COL[9977] = 1'b1;
assign COL[9978] = 1'b1;
assign COL[9979] = 1'b1;
assign COL[9980] = 1'b1;
assign COL[9981] = 1'b1;
assign COL[9982] = 1'b0;
assign COL[9983] = 1'b0;
assign COL[9984] = 1'b0;
assign COL[9985] = 1'b0;
assign COL[9986] = 1'b0;
assign COL[9987] = 1'b0;
assign COL[9988] = 1'b0;
assign COL[9989] = 1'b0;
assign COL[9990] = 1'b1;
assign COL[9991] = 1'b1;
assign COL[9992] = 1'b1;
assign COL[9993] = 1'b1;
assign COL[9994] = 1'b1;
assign COL[9995] = 1'b1;
assign COL[9996] = 1'b1;
assign COL[9997] = 1'b1;
assign COL[9998] = 1'b1;
assign COL[9999] = 1'b1;
assign COL[10000] = 1'b1;
assign COL[10001] = 1'b1;
assign COL[10002] = 1'b1;
assign COL[10003] = 1'b1;
assign COL[10004] = 1'b1;
assign COL[10005] = 1'b1;
assign COL[10006] = 1'b1;
assign COL[10007] = 1'b1;
assign COL[10008] = 1'b1;
assign COL[10009] = 1'b1;
assign COL[10010] = 1'b1;
assign COL[10011] = 1'b1;
assign COL[10012] = 1'b1;
assign COL[10013] = 1'b1;
assign COL[10014] = 1'b1;
assign COL[10015] = 1'b0;
assign COL[10016] = 1'b0;
assign COL[10017] = 1'b0;
assign COL[10018] = 1'b0;
assign COL[10019] = 1'b0;
assign COL[10020] = 1'b0;
assign COL[10021] = 1'b0;
assign COL[10022] = 1'b0;
assign COL[10023] = 1'b0;
assign COL[10024] = 1'b0;
assign COL[10025] = 1'b0;
assign COL[10026] = 1'b0;
assign COL[10027] = 1'b0;
assign COL[10028] = 1'b0;
assign COL[10029] = 1'b0;
assign COL[10030] = 1'b0;
assign COL[10031] = 1'b0;
assign COL[10032] = 1'b0;
assign COL[10033] = 1'b0;
assign COL[10034] = 1'b0;
assign COL[10035] = 1'b0;
assign COL[10036] = 1'b0;
assign COL[10037] = 1'b0;
assign COL[10038] = 1'b0;
assign COL[10039] = 1'b0;
assign COL[10040] = 1'b0;
assign COL[10041] = 1'b0;
assign COL[10042] = 1'b0;
assign COL[10043] = 1'b0;
assign COL[10044] = 1'b0;
assign COL[10045] = 1'b0;
assign COL[10046] = 1'b0;
assign COL[10047] = 1'b0;
assign COL[10048] = 1'b0;
assign COL[10049] = 1'b0;
assign COL[10050] = 1'b0;
assign COL[10051] = 1'b0;
assign COL[10052] = 1'b0;
assign COL[10053] = 1'b0;
assign COL[10054] = 1'b0;
assign COL[10055] = 1'b0;
assign COL[10056] = 1'b0;
assign COL[10057] = 1'b0;
assign COL[10058] = 1'b0;
assign COL[10059] = 1'b0;
assign COL[10060] = 1'b0;
assign COL[10061] = 1'b0;
assign COL[10062] = 1'b0;
assign COL[10063] = 1'b0;
assign COL[10064] = 1'b0;
assign COL[10065] = 1'b0;
assign COL[10066] = 1'b0;
assign COL[10067] = 1'b0;
assign COL[10068] = 1'b0;
assign COL[10069] = 1'b0;
assign COL[10070] = 1'b0;
assign COL[10071] = 1'b0;
assign COL[10072] = 1'b0;
assign COL[10073] = 1'b0;
assign COL[10074] = 1'b0;
assign COL[10075] = 1'b0;
assign COL[10076] = 1'b0;
assign COL[10077] = 1'b0;
assign COL[10078] = 1'b0;
assign COL[10079] = 1'b0;
assign COL[10080] = 1'b0;
assign COL[10081] = 1'b1;
assign COL[10082] = 1'b1;
assign COL[10083] = 1'b1;
assign COL[10084] = 1'b1;
assign COL[10085] = 1'b1;
assign COL[10086] = 1'b1;
assign COL[10087] = 1'b1;
assign COL[10088] = 1'b1;
assign COL[10089] = 1'b1;
assign COL[10090] = 1'b1;
assign COL[10091] = 1'b1;
assign COL[10092] = 1'b1;
assign COL[10093] = 1'b1;
assign COL[10094] = 1'b1;
assign COL[10095] = 1'b0;
assign COL[10096] = 1'b0;
assign COL[10097] = 1'b0;
assign COL[10098] = 1'b0;
assign COL[10099] = 1'b0;
assign COL[10100] = 1'b0;
assign COL[10101] = 1'b0;
assign COL[10102] = 1'b0;
assign COL[10103] = 1'b0;
assign COL[10104] = 1'b0;
assign COL[10105] = 1'b0;
assign COL[10106] = 1'b0;
assign COL[10107] = 1'b0;
assign COL[10108] = 1'b0;
assign COL[10109] = 1'b1;
assign COL[10110] = 1'b1;
assign COL[10111] = 1'b1;
assign COL[10112] = 1'b1;
assign COL[10113] = 1'b0;
assign COL[10114] = 1'b0;
assign COL[10115] = 1'b0;
assign COL[10116] = 1'b0;
assign COL[10117] = 1'b0;
assign COL[10118] = 1'b0;
assign COL[10119] = 1'b0;
assign COL[10120] = 1'b0;
assign COL[10121] = 1'b0;
assign COL[10122] = 1'b0;
assign COL[10123] = 1'b0;
assign COL[10124] = 1'b0;
assign COL[10125] = 1'b1;
assign COL[10126] = 1'b1;
assign COL[10127] = 1'b1;
assign COL[10128] = 1'b1;
assign COL[10129] = 1'b1;
assign COL[10130] = 1'b1;
assign COL[10131] = 1'b1;
assign COL[10132] = 1'b1;
assign COL[10133] = 1'b1;
assign COL[10134] = 1'b1;
assign COL[10135] = 1'b1;
assign COL[10136] = 1'b1;
assign COL[10137] = 1'b1;
assign COL[10138] = 1'b1;
assign COL[10139] = 1'b1;
assign COL[10140] = 1'b1;
assign COL[10141] = 1'b1;
assign COL[10142] = 1'b0;
assign COL[10143] = 1'b0;
assign COL[10144] = 1'b0;
assign COL[10145] = 1'b0;
assign COL[10146] = 1'b0;
assign COL[10147] = 1'b0;
assign COL[10148] = 1'b0;
assign COL[10149] = 1'b0;
assign COL[10150] = 1'b1;
assign COL[10151] = 1'b1;
assign COL[10152] = 1'b1;
assign COL[10153] = 1'b1;
assign COL[10154] = 1'b1;
assign COL[10155] = 1'b1;
assign COL[10156] = 1'b1;
assign COL[10157] = 1'b1;
assign COL[10158] = 1'b1;
assign COL[10159] = 1'b1;
assign COL[10160] = 1'b1;
assign COL[10161] = 1'b1;
assign COL[10162] = 1'b1;
assign COL[10163] = 1'b1;
assign COL[10164] = 1'b1;
assign COL[10165] = 1'b1;
assign COL[10166] = 1'b1;
assign COL[10167] = 1'b1;
assign COL[10168] = 1'b1;
assign COL[10169] = 1'b1;
assign COL[10170] = 1'b1;
assign COL[10171] = 1'b1;
assign COL[10172] = 1'b1;
assign COL[10173] = 1'b1;
assign COL[10174] = 1'b1;
assign COL[10175] = 1'b0;
assign COL[10176] = 1'b0;
assign COL[10177] = 1'b0;
assign COL[10178] = 1'b0;
assign COL[10179] = 1'b0;
assign COL[10180] = 1'b0;
assign COL[10181] = 1'b0;
assign COL[10182] = 1'b0;
assign COL[10183] = 1'b0;
assign COL[10184] = 1'b0;
assign COL[10185] = 1'b0;
assign COL[10186] = 1'b0;
assign COL[10187] = 1'b0;
assign COL[10188] = 1'b0;
assign COL[10189] = 1'b0;
assign COL[10190] = 1'b0;
assign COL[10191] = 1'b0;
assign COL[10192] = 1'b0;
assign COL[10193] = 1'b0;
assign COL[10194] = 1'b0;
assign COL[10195] = 1'b0;
assign COL[10196] = 1'b0;
assign COL[10197] = 1'b0;
assign COL[10198] = 1'b0;
assign COL[10199] = 1'b0;
assign COL[10200] = 1'b0;
assign COL[10201] = 1'b0;
assign COL[10202] = 1'b0;
assign COL[10203] = 1'b0;
assign COL[10204] = 1'b0;
assign COL[10205] = 1'b0;
assign COL[10206] = 1'b0;
assign COL[10207] = 1'b0;
assign COL[10208] = 1'b0;
assign COL[10209] = 1'b0;
assign COL[10210] = 1'b0;
assign COL[10211] = 1'b0;
assign COL[10212] = 1'b0;
assign COL[10213] = 1'b0;
assign COL[10214] = 1'b0;
assign COL[10215] = 1'b0;
assign COL[10216] = 1'b0;
assign COL[10217] = 1'b0;
assign COL[10218] = 1'b0;
assign COL[10219] = 1'b0;
assign COL[10220] = 1'b0;
assign COL[10221] = 1'b0;
assign COL[10222] = 1'b0;
assign COL[10223] = 1'b0;
assign COL[10224] = 1'b0;
assign COL[10225] = 1'b0;
assign COL[10226] = 1'b0;
assign COL[10227] = 1'b0;
assign COL[10228] = 1'b0;
assign COL[10229] = 1'b0;
assign COL[10230] = 1'b0;
assign COL[10231] = 1'b0;
assign COL[10232] = 1'b0;
assign COL[10233] = 1'b0;
assign COL[10234] = 1'b0;
assign COL[10235] = 1'b0;
assign COL[10236] = 1'b0;
assign COL[10237] = 1'b0;
assign COL[10238] = 1'b0;
assign COL[10239] = 1'b0;
assign COL[10240] = 1'b0;
assign COL[10241] = 1'b1;
assign COL[10242] = 1'b1;
assign COL[10243] = 1'b1;
assign COL[10244] = 1'b1;
assign COL[10245] = 1'b1;
assign COL[10246] = 1'b1;
assign COL[10247] = 1'b1;
assign COL[10248] = 1'b1;
assign COL[10249] = 1'b1;
assign COL[10250] = 1'b1;
assign COL[10251] = 1'b1;
assign COL[10252] = 1'b1;
assign COL[10253] = 1'b1;
assign COL[10254] = 1'b1;
assign COL[10255] = 1'b0;
assign COL[10256] = 1'b0;
assign COL[10257] = 1'b0;
assign COL[10258] = 1'b0;
assign COL[10259] = 1'b0;
assign COL[10260] = 1'b0;
assign COL[10261] = 1'b0;
assign COL[10262] = 1'b0;
assign COL[10263] = 1'b0;
assign COL[10264] = 1'b0;
assign COL[10265] = 1'b0;
assign COL[10266] = 1'b0;
assign COL[10267] = 1'b0;
assign COL[10268] = 1'b0;
assign COL[10269] = 1'b1;
assign COL[10270] = 1'b1;
assign COL[10271] = 1'b1;
assign COL[10272] = 1'b1;
assign COL[10273] = 1'b0;
assign COL[10274] = 1'b0;
assign COL[10275] = 1'b0;
assign COL[10276] = 1'b0;
assign COL[10277] = 1'b0;
assign COL[10278] = 1'b0;
assign COL[10279] = 1'b0;
assign COL[10280] = 1'b0;
assign COL[10281] = 1'b0;
assign COL[10282] = 1'b0;
assign COL[10283] = 1'b0;
assign COL[10284] = 1'b0;
assign COL[10285] = 1'b1;
assign COL[10286] = 1'b1;
assign COL[10287] = 1'b1;
assign COL[10288] = 1'b1;
assign COL[10289] = 1'b1;
assign COL[10290] = 1'b1;
assign COL[10291] = 1'b1;
assign COL[10292] = 1'b1;
assign COL[10293] = 1'b1;
assign COL[10294] = 1'b1;
assign COL[10295] = 1'b1;
assign COL[10296] = 1'b1;
assign COL[10297] = 1'b1;
assign COL[10298] = 1'b1;
assign COL[10299] = 1'b1;
assign COL[10300] = 1'b1;
assign COL[10301] = 1'b1;
assign COL[10302] = 1'b0;
assign COL[10303] = 1'b0;
assign COL[10304] = 1'b0;
assign COL[10305] = 1'b0;
assign COL[10306] = 1'b0;
assign COL[10307] = 1'b0;
assign COL[10308] = 1'b0;
assign COL[10309] = 1'b0;
assign COL[10310] = 1'b1;
assign COL[10311] = 1'b1;
assign COL[10312] = 1'b1;
assign COL[10313] = 1'b1;
assign COL[10314] = 1'b1;
assign COL[10315] = 1'b1;
assign COL[10316] = 1'b1;
assign COL[10317] = 1'b1;
assign COL[10318] = 1'b1;
assign COL[10319] = 1'b1;
assign COL[10320] = 1'b1;
assign COL[10321] = 1'b1;
assign COL[10322] = 1'b1;
assign COL[10323] = 1'b1;
assign COL[10324] = 1'b1;
assign COL[10325] = 1'b1;
assign COL[10326] = 1'b1;
assign COL[10327] = 1'b1;
assign COL[10328] = 1'b1;
assign COL[10329] = 1'b1;
assign COL[10330] = 1'b1;
assign COL[10331] = 1'b1;
assign COL[10332] = 1'b1;
assign COL[10333] = 1'b1;
assign COL[10334] = 1'b1;
assign COL[10335] = 1'b0;
assign COL[10336] = 1'b0;
assign COL[10337] = 1'b0;
assign COL[10338] = 1'b0;
assign COL[10339] = 1'b0;
assign COL[10340] = 1'b0;
assign COL[10341] = 1'b0;
assign COL[10342] = 1'b0;
assign COL[10343] = 1'b0;
assign COL[10344] = 1'b0;
assign COL[10345] = 1'b0;
assign COL[10346] = 1'b0;
assign COL[10347] = 1'b0;
assign COL[10348] = 1'b0;
assign COL[10349] = 1'b0;
assign COL[10350] = 1'b0;
assign COL[10351] = 1'b0;
assign COL[10352] = 1'b0;
assign COL[10353] = 1'b0;
assign COL[10354] = 1'b0;
assign COL[10355] = 1'b0;
assign COL[10356] = 1'b0;
assign COL[10357] = 1'b0;
assign COL[10358] = 1'b0;
assign COL[10359] = 1'b0;
assign COL[10360] = 1'b0;
assign COL[10361] = 1'b0;
assign COL[10362] = 1'b0;
assign COL[10363] = 1'b0;
assign COL[10364] = 1'b0;
assign COL[10365] = 1'b0;
assign COL[10366] = 1'b0;
assign COL[10367] = 1'b0;
assign COL[10368] = 1'b0;
assign COL[10369] = 1'b0;
assign COL[10370] = 1'b0;
assign COL[10371] = 1'b0;
assign COL[10372] = 1'b0;
assign COL[10373] = 1'b0;
assign COL[10374] = 1'b0;
assign COL[10375] = 1'b0;
assign COL[10376] = 1'b0;
assign COL[10377] = 1'b0;
assign COL[10378] = 1'b0;
assign COL[10379] = 1'b0;
assign COL[10380] = 1'b0;
assign COL[10381] = 1'b0;
assign COL[10382] = 1'b0;
assign COL[10383] = 1'b0;
assign COL[10384] = 1'b0;
assign COL[10385] = 1'b0;
assign COL[10386] = 1'b0;
assign COL[10387] = 1'b0;
assign COL[10388] = 1'b0;
assign COL[10389] = 1'b0;
assign COL[10390] = 1'b0;
assign COL[10391] = 1'b0;
assign COL[10392] = 1'b0;
assign COL[10393] = 1'b0;
assign COL[10394] = 1'b0;
assign COL[10395] = 1'b0;
assign COL[10396] = 1'b0;
assign COL[10397] = 1'b0;
assign COL[10398] = 1'b0;
assign COL[10399] = 1'b0;
assign COL[10400] = 1'b0;
assign COL[10401] = 1'b1;
assign COL[10402] = 1'b1;
assign COL[10403] = 1'b1;
assign COL[10404] = 1'b1;
assign COL[10405] = 1'b1;
assign COL[10406] = 1'b1;
assign COL[10407] = 1'b1;
assign COL[10408] = 1'b1;
assign COL[10409] = 1'b1;
assign COL[10410] = 1'b1;
assign COL[10411] = 1'b1;
assign COL[10412] = 1'b1;
assign COL[10413] = 1'b1;
assign COL[10414] = 1'b1;
assign COL[10415] = 1'b0;
assign COL[10416] = 1'b0;
assign COL[10417] = 1'b0;
assign COL[10418] = 1'b0;
assign COL[10419] = 1'b0;
assign COL[10420] = 1'b0;
assign COL[10421] = 1'b0;
assign COL[10422] = 1'b0;
assign COL[10423] = 1'b0;
assign COL[10424] = 1'b0;
assign COL[10425] = 1'b0;
assign COL[10426] = 1'b0;
assign COL[10427] = 1'b0;
assign COL[10428] = 1'b0;
assign COL[10429] = 1'b1;
assign COL[10430] = 1'b1;
assign COL[10431] = 1'b1;
assign COL[10432] = 1'b1;
assign COL[10433] = 1'b0;
assign COL[10434] = 1'b0;
assign COL[10435] = 1'b0;
assign COL[10436] = 1'b0;
assign COL[10437] = 1'b0;
assign COL[10438] = 1'b0;
assign COL[10439] = 1'b0;
assign COL[10440] = 1'b0;
assign COL[10441] = 1'b0;
assign COL[10442] = 1'b0;
assign COL[10443] = 1'b0;
assign COL[10444] = 1'b0;
assign COL[10445] = 1'b1;
assign COL[10446] = 1'b1;
assign COL[10447] = 1'b1;
assign COL[10448] = 1'b1;
assign COL[10449] = 1'b1;
assign COL[10450] = 1'b1;
assign COL[10451] = 1'b1;
assign COL[10452] = 1'b1;
assign COL[10453] = 1'b1;
assign COL[10454] = 1'b1;
assign COL[10455] = 1'b1;
assign COL[10456] = 1'b1;
assign COL[10457] = 1'b1;
assign COL[10458] = 1'b1;
assign COL[10459] = 1'b1;
assign COL[10460] = 1'b1;
assign COL[10461] = 1'b1;
assign COL[10462] = 1'b0;
assign COL[10463] = 1'b0;
assign COL[10464] = 1'b0;
assign COL[10465] = 1'b0;
assign COL[10466] = 1'b0;
assign COL[10467] = 1'b0;
assign COL[10468] = 1'b0;
assign COL[10469] = 1'b0;
assign COL[10470] = 1'b1;
assign COL[10471] = 1'b1;
assign COL[10472] = 1'b1;
assign COL[10473] = 1'b1;
assign COL[10474] = 1'b1;
assign COL[10475] = 1'b1;
assign COL[10476] = 1'b1;
assign COL[10477] = 1'b1;
assign COL[10478] = 1'b1;
assign COL[10479] = 1'b1;
assign COL[10480] = 1'b1;
assign COL[10481] = 1'b1;
assign COL[10482] = 1'b1;
assign COL[10483] = 1'b1;
assign COL[10484] = 1'b1;
assign COL[10485] = 1'b1;
assign COL[10486] = 1'b1;
assign COL[10487] = 1'b1;
assign COL[10488] = 1'b1;
assign COL[10489] = 1'b1;
assign COL[10490] = 1'b1;
assign COL[10491] = 1'b1;
assign COL[10492] = 1'b1;
assign COL[10493] = 1'b1;
assign COL[10494] = 1'b1;
assign COL[10495] = 1'b0;
assign COL[10496] = 1'b0;
assign COL[10497] = 1'b0;
assign COL[10498] = 1'b0;
assign COL[10499] = 1'b0;
assign COL[10500] = 1'b0;
assign COL[10501] = 1'b0;
assign COL[10502] = 1'b0;
assign COL[10503] = 1'b0;
assign COL[10504] = 1'b0;
assign COL[10505] = 1'b0;
assign COL[10506] = 1'b0;
assign COL[10507] = 1'b0;
assign COL[10508] = 1'b0;
assign COL[10509] = 1'b0;
assign COL[10510] = 1'b0;
assign COL[10511] = 1'b0;
assign COL[10512] = 1'b0;
assign COL[10513] = 1'b0;
assign COL[10514] = 1'b0;
assign COL[10515] = 1'b0;
assign COL[10516] = 1'b0;
assign COL[10517] = 1'b0;
assign COL[10518] = 1'b0;
assign COL[10519] = 1'b0;
assign COL[10520] = 1'b0;
assign COL[10521] = 1'b0;
assign COL[10522] = 1'b0;
assign COL[10523] = 1'b0;
assign COL[10524] = 1'b0;
assign COL[10525] = 1'b0;
assign COL[10526] = 1'b0;
assign COL[10527] = 1'b0;
assign COL[10528] = 1'b0;
assign COL[10529] = 1'b0;
assign COL[10530] = 1'b0;
assign COL[10531] = 1'b0;
assign COL[10532] = 1'b0;
assign COL[10533] = 1'b0;
assign COL[10534] = 1'b0;
assign COL[10535] = 1'b0;
assign COL[10536] = 1'b0;
assign COL[10537] = 1'b0;
assign COL[10538] = 1'b0;
assign COL[10539] = 1'b0;
assign COL[10540] = 1'b0;
assign COL[10541] = 1'b0;
assign COL[10542] = 1'b0;
assign COL[10543] = 1'b0;
assign COL[10544] = 1'b0;
assign COL[10545] = 1'b0;
assign COL[10546] = 1'b0;
assign COL[10547] = 1'b0;
assign COL[10548] = 1'b0;
assign COL[10549] = 1'b0;
assign COL[10550] = 1'b0;
assign COL[10551] = 1'b0;
assign COL[10552] = 1'b0;
assign COL[10553] = 1'b0;
assign COL[10554] = 1'b0;
assign COL[10555] = 1'b0;
assign COL[10556] = 1'b0;
assign COL[10557] = 1'b0;
assign COL[10558] = 1'b0;
assign COL[10559] = 1'b0;
assign COL[10560] = 1'b0;
assign COL[10561] = 1'b1;
assign COL[10562] = 1'b1;
assign COL[10563] = 1'b1;
assign COL[10564] = 1'b1;
assign COL[10565] = 1'b1;
assign COL[10566] = 1'b1;
assign COL[10567] = 1'b1;
assign COL[10568] = 1'b1;
assign COL[10569] = 1'b1;
assign COL[10570] = 1'b1;
assign COL[10571] = 1'b1;
assign COL[10572] = 1'b1;
assign COL[10573] = 1'b1;
assign COL[10574] = 1'b1;
assign COL[10575] = 1'b0;
assign COL[10576] = 1'b0;
assign COL[10577] = 1'b0;
assign COL[10578] = 1'b0;
assign COL[10579] = 1'b0;
assign COL[10580] = 1'b0;
assign COL[10581] = 1'b0;
assign COL[10582] = 1'b0;
assign COL[10583] = 1'b0;
assign COL[10584] = 1'b0;
assign COL[10585] = 1'b0;
assign COL[10586] = 1'b0;
assign COL[10587] = 1'b0;
assign COL[10588] = 1'b0;
assign COL[10589] = 1'b1;
assign COL[10590] = 1'b1;
assign COL[10591] = 1'b1;
assign COL[10592] = 1'b1;
assign COL[10593] = 1'b0;
assign COL[10594] = 1'b0;
assign COL[10595] = 1'b0;
assign COL[10596] = 1'b0;
assign COL[10597] = 1'b0;
assign COL[10598] = 1'b0;
assign COL[10599] = 1'b0;
assign COL[10600] = 1'b0;
assign COL[10601] = 1'b0;
assign COL[10602] = 1'b0;
assign COL[10603] = 1'b0;
assign COL[10604] = 1'b0;
assign COL[10605] = 1'b1;
assign COL[10606] = 1'b1;
assign COL[10607] = 1'b1;
assign COL[10608] = 1'b1;
assign COL[10609] = 1'b0;
assign COL[10610] = 1'b0;
assign COL[10611] = 1'b0;
assign COL[10612] = 1'b0;
assign COL[10613] = 1'b0;
assign COL[10614] = 1'b0;
assign COL[10615] = 1'b0;
assign COL[10616] = 1'b0;
assign COL[10617] = 1'b0;
assign COL[10618] = 1'b0;
assign COL[10619] = 1'b0;
assign COL[10620] = 1'b0;
assign COL[10621] = 1'b0;
assign COL[10622] = 1'b0;
assign COL[10623] = 1'b0;
assign COL[10624] = 1'b0;
assign COL[10625] = 1'b0;
assign COL[10626] = 1'b0;
assign COL[10627] = 1'b0;
assign COL[10628] = 1'b0;
assign COL[10629] = 1'b0;
assign COL[10630] = 1'b0;
assign COL[10631] = 1'b0;
assign COL[10632] = 1'b0;
assign COL[10633] = 1'b0;
assign COL[10634] = 1'b0;
assign COL[10635] = 1'b0;
assign COL[10636] = 1'b0;
assign COL[10637] = 1'b0;
assign COL[10638] = 1'b0;
assign COL[10639] = 1'b0;
assign COL[10640] = 1'b0;
assign COL[10641] = 1'b0;
assign COL[10642] = 1'b0;
assign COL[10643] = 1'b0;
assign COL[10644] = 1'b0;
assign COL[10645] = 1'b0;
assign COL[10646] = 1'b0;
assign COL[10647] = 1'b0;
assign COL[10648] = 1'b0;
assign COL[10649] = 1'b0;
assign COL[10650] = 1'b1;
assign COL[10651] = 1'b1;
assign COL[10652] = 1'b1;
assign COL[10653] = 1'b1;
assign COL[10654] = 1'b1;
assign COL[10655] = 1'b0;
assign COL[10656] = 1'b0;
assign COL[10657] = 1'b0;
assign COL[10658] = 1'b0;
assign COL[10659] = 1'b0;
assign COL[10660] = 1'b0;
assign COL[10661] = 1'b0;
assign COL[10662] = 1'b0;
assign COL[10663] = 1'b0;
assign COL[10664] = 1'b0;
assign COL[10665] = 1'b0;
assign COL[10666] = 1'b0;
assign COL[10667] = 1'b0;
assign COL[10668] = 1'b0;
assign COL[10669] = 1'b0;
assign COL[10670] = 1'b0;
assign COL[10671] = 1'b0;
assign COL[10672] = 1'b0;
assign COL[10673] = 1'b0;
assign COL[10674] = 1'b0;
assign COL[10675] = 1'b0;
assign COL[10676] = 1'b0;
assign COL[10677] = 1'b0;
assign COL[10678] = 1'b0;
assign COL[10679] = 1'b0;
assign COL[10680] = 1'b0;
assign COL[10681] = 1'b0;
assign COL[10682] = 1'b0;
assign COL[10683] = 1'b0;
assign COL[10684] = 1'b0;
assign COL[10685] = 1'b0;
assign COL[10686] = 1'b0;
assign COL[10687] = 1'b0;
assign COL[10688] = 1'b0;
assign COL[10689] = 1'b0;
assign COL[10690] = 1'b0;
assign COL[10691] = 1'b0;
assign COL[10692] = 1'b0;
assign COL[10693] = 1'b0;
assign COL[10694] = 1'b0;
assign COL[10695] = 1'b0;
assign COL[10696] = 1'b0;
assign COL[10697] = 1'b0;
assign COL[10698] = 1'b0;
assign COL[10699] = 1'b0;
assign COL[10700] = 1'b0;
assign COL[10701] = 1'b0;
assign COL[10702] = 1'b0;
assign COL[10703] = 1'b0;
assign COL[10704] = 1'b0;
assign COL[10705] = 1'b0;
assign COL[10706] = 1'b0;
assign COL[10707] = 1'b0;
assign COL[10708] = 1'b0;
assign COL[10709] = 1'b0;
assign COL[10710] = 1'b0;
assign COL[10711] = 1'b0;
assign COL[10712] = 1'b0;
assign COL[10713] = 1'b0;
assign COL[10714] = 1'b0;
assign COL[10715] = 1'b0;
assign COL[10716] = 1'b0;
assign COL[10717] = 1'b0;
assign COL[10718] = 1'b0;
assign COL[10719] = 1'b0;
assign COL[10720] = 1'b0;
assign COL[10721] = 1'b1;
assign COL[10722] = 1'b1;
assign COL[10723] = 1'b1;
assign COL[10724] = 1'b1;
assign COL[10725] = 1'b0;
assign COL[10726] = 1'b0;
assign COL[10727] = 1'b0;
assign COL[10728] = 1'b0;
assign COL[10729] = 1'b0;
assign COL[10730] = 1'b0;
assign COL[10731] = 1'b0;
assign COL[10732] = 1'b0;
assign COL[10733] = 1'b0;
assign COL[10734] = 1'b0;
assign COL[10735] = 1'b0;
assign COL[10736] = 1'b0;
assign COL[10737] = 1'b0;
assign COL[10738] = 1'b0;
assign COL[10739] = 1'b0;
assign COL[10740] = 1'b0;
assign COL[10741] = 1'b0;
assign COL[10742] = 1'b0;
assign COL[10743] = 1'b0;
assign COL[10744] = 1'b0;
assign COL[10745] = 1'b0;
assign COL[10746] = 1'b0;
assign COL[10747] = 1'b0;
assign COL[10748] = 1'b0;
assign COL[10749] = 1'b1;
assign COL[10750] = 1'b1;
assign COL[10751] = 1'b1;
assign COL[10752] = 1'b1;
assign COL[10753] = 1'b0;
assign COL[10754] = 1'b0;
assign COL[10755] = 1'b0;
assign COL[10756] = 1'b0;
assign COL[10757] = 1'b0;
assign COL[10758] = 1'b0;
assign COL[10759] = 1'b0;
assign COL[10760] = 1'b0;
assign COL[10761] = 1'b0;
assign COL[10762] = 1'b0;
assign COL[10763] = 1'b0;
assign COL[10764] = 1'b0;
assign COL[10765] = 1'b1;
assign COL[10766] = 1'b1;
assign COL[10767] = 1'b1;
assign COL[10768] = 1'b1;
assign COL[10769] = 1'b0;
assign COL[10770] = 1'b0;
assign COL[10771] = 1'b0;
assign COL[10772] = 1'b0;
assign COL[10773] = 1'b0;
assign COL[10774] = 1'b0;
assign COL[10775] = 1'b0;
assign COL[10776] = 1'b0;
assign COL[10777] = 1'b0;
assign COL[10778] = 1'b0;
assign COL[10779] = 1'b0;
assign COL[10780] = 1'b0;
assign COL[10781] = 1'b0;
assign COL[10782] = 1'b0;
assign COL[10783] = 1'b0;
assign COL[10784] = 1'b0;
assign COL[10785] = 1'b0;
assign COL[10786] = 1'b0;
assign COL[10787] = 1'b0;
assign COL[10788] = 1'b0;
assign COL[10789] = 1'b0;
assign COL[10790] = 1'b0;
assign COL[10791] = 1'b0;
assign COL[10792] = 1'b0;
assign COL[10793] = 1'b0;
assign COL[10794] = 1'b0;
assign COL[10795] = 1'b0;
assign COL[10796] = 1'b0;
assign COL[10797] = 1'b0;
assign COL[10798] = 1'b0;
assign COL[10799] = 1'b0;
assign COL[10800] = 1'b0;
assign COL[10801] = 1'b0;
assign COL[10802] = 1'b0;
assign COL[10803] = 1'b0;
assign COL[10804] = 1'b0;
assign COL[10805] = 1'b0;
assign COL[10806] = 1'b0;
assign COL[10807] = 1'b0;
assign COL[10808] = 1'b0;
assign COL[10809] = 1'b0;
assign COL[10810] = 1'b1;
assign COL[10811] = 1'b1;
assign COL[10812] = 1'b1;
assign COL[10813] = 1'b1;
assign COL[10814] = 1'b1;
assign COL[10815] = 1'b0;
assign COL[10816] = 1'b0;
assign COL[10817] = 1'b0;
assign COL[10818] = 1'b0;
assign COL[10819] = 1'b0;
assign COL[10820] = 1'b0;
assign COL[10821] = 1'b0;
assign COL[10822] = 1'b0;
assign COL[10823] = 1'b0;
assign COL[10824] = 1'b0;
assign COL[10825] = 1'b0;
assign COL[10826] = 1'b0;
assign COL[10827] = 1'b0;
assign COL[10828] = 1'b0;
assign COL[10829] = 1'b0;
assign COL[10830] = 1'b0;
assign COL[10831] = 1'b0;
assign COL[10832] = 1'b0;
assign COL[10833] = 1'b0;
assign COL[10834] = 1'b0;
assign COL[10835] = 1'b0;
assign COL[10836] = 1'b0;
assign COL[10837] = 1'b0;
assign COL[10838] = 1'b0;
assign COL[10839] = 1'b0;
assign COL[10840] = 1'b0;
assign COL[10841] = 1'b0;
assign COL[10842] = 1'b0;
assign COL[10843] = 1'b0;
assign COL[10844] = 1'b0;
assign COL[10845] = 1'b0;
assign COL[10846] = 1'b0;
assign COL[10847] = 1'b0;
assign COL[10848] = 1'b0;
assign COL[10849] = 1'b0;
assign COL[10850] = 1'b0;
assign COL[10851] = 1'b0;
assign COL[10852] = 1'b0;
assign COL[10853] = 1'b0;
assign COL[10854] = 1'b0;
assign COL[10855] = 1'b0;
assign COL[10856] = 1'b0;
assign COL[10857] = 1'b0;
assign COL[10858] = 1'b0;
assign COL[10859] = 1'b0;
assign COL[10860] = 1'b0;
assign COL[10861] = 1'b0;
assign COL[10862] = 1'b0;
assign COL[10863] = 1'b0;
assign COL[10864] = 1'b0;
assign COL[10865] = 1'b0;
assign COL[10866] = 1'b0;
assign COL[10867] = 1'b0;
assign COL[10868] = 1'b0;
assign COL[10869] = 1'b0;
assign COL[10870] = 1'b0;
assign COL[10871] = 1'b0;
assign COL[10872] = 1'b0;
assign COL[10873] = 1'b0;
assign COL[10874] = 1'b0;
assign COL[10875] = 1'b0;
assign COL[10876] = 1'b0;
assign COL[10877] = 1'b0;
assign COL[10878] = 1'b0;
assign COL[10879] = 1'b0;
assign COL[10880] = 1'b0;
assign COL[10881] = 1'b1;
assign COL[10882] = 1'b1;
assign COL[10883] = 1'b1;
assign COL[10884] = 1'b1;
assign COL[10885] = 1'b0;
assign COL[10886] = 1'b0;
assign COL[10887] = 1'b0;
assign COL[10888] = 1'b0;
assign COL[10889] = 1'b0;
assign COL[10890] = 1'b0;
assign COL[10891] = 1'b0;
assign COL[10892] = 1'b0;
assign COL[10893] = 1'b0;
assign COL[10894] = 1'b0;
assign COL[10895] = 1'b0;
assign COL[10896] = 1'b0;
assign COL[10897] = 1'b0;
assign COL[10898] = 1'b0;
assign COL[10899] = 1'b0;
assign COL[10900] = 1'b0;
assign COL[10901] = 1'b0;
assign COL[10902] = 1'b0;
assign COL[10903] = 1'b0;
assign COL[10904] = 1'b0;
assign COL[10905] = 1'b0;
assign COL[10906] = 1'b0;
assign COL[10907] = 1'b0;
assign COL[10908] = 1'b0;
assign COL[10909] = 1'b1;
assign COL[10910] = 1'b1;
assign COL[10911] = 1'b1;
assign COL[10912] = 1'b1;
assign COL[10913] = 1'b0;
assign COL[10914] = 1'b0;
assign COL[10915] = 1'b0;
assign COL[10916] = 1'b0;
assign COL[10917] = 1'b0;
assign COL[10918] = 1'b0;
assign COL[10919] = 1'b0;
assign COL[10920] = 1'b0;
assign COL[10921] = 1'b0;
assign COL[10922] = 1'b0;
assign COL[10923] = 1'b0;
assign COL[10924] = 1'b0;
assign COL[10925] = 1'b1;
assign COL[10926] = 1'b1;
assign COL[10927] = 1'b1;
assign COL[10928] = 1'b1;
assign COL[10929] = 1'b0;
assign COL[10930] = 1'b0;
assign COL[10931] = 1'b0;
assign COL[10932] = 1'b0;
assign COL[10933] = 1'b0;
assign COL[10934] = 1'b0;
assign COL[10935] = 1'b0;
assign COL[10936] = 1'b0;
assign COL[10937] = 1'b0;
assign COL[10938] = 1'b0;
assign COL[10939] = 1'b0;
assign COL[10940] = 1'b0;
assign COL[10941] = 1'b0;
assign COL[10942] = 1'b0;
assign COL[10943] = 1'b0;
assign COL[10944] = 1'b0;
assign COL[10945] = 1'b0;
assign COL[10946] = 1'b0;
assign COL[10947] = 1'b0;
assign COL[10948] = 1'b0;
assign COL[10949] = 1'b0;
assign COL[10950] = 1'b0;
assign COL[10951] = 1'b0;
assign COL[10952] = 1'b0;
assign COL[10953] = 1'b0;
assign COL[10954] = 1'b0;
assign COL[10955] = 1'b0;
assign COL[10956] = 1'b0;
assign COL[10957] = 1'b0;
assign COL[10958] = 1'b0;
assign COL[10959] = 1'b0;
assign COL[10960] = 1'b0;
assign COL[10961] = 1'b0;
assign COL[10962] = 1'b0;
assign COL[10963] = 1'b0;
assign COL[10964] = 1'b0;
assign COL[10965] = 1'b0;
assign COL[10966] = 1'b0;
assign COL[10967] = 1'b0;
assign COL[10968] = 1'b0;
assign COL[10969] = 1'b0;
assign COL[10970] = 1'b1;
assign COL[10971] = 1'b1;
assign COL[10972] = 1'b1;
assign COL[10973] = 1'b1;
assign COL[10974] = 1'b1;
assign COL[10975] = 1'b0;
assign COL[10976] = 1'b0;
assign COL[10977] = 1'b0;
assign COL[10978] = 1'b0;
assign COL[10979] = 1'b0;
assign COL[10980] = 1'b0;
assign COL[10981] = 1'b0;
assign COL[10982] = 1'b0;
assign COL[10983] = 1'b0;
assign COL[10984] = 1'b0;
assign COL[10985] = 1'b0;
assign COL[10986] = 1'b0;
assign COL[10987] = 1'b0;
assign COL[10988] = 1'b0;
assign COL[10989] = 1'b0;
assign COL[10990] = 1'b0;
assign COL[10991] = 1'b0;
assign COL[10992] = 1'b0;
assign COL[10993] = 1'b0;
assign COL[10994] = 1'b0;
assign COL[10995] = 1'b0;
assign COL[10996] = 1'b0;
assign COL[10997] = 1'b0;
assign COL[10998] = 1'b0;
assign COL[10999] = 1'b0;
assign COL[11000] = 1'b0;
assign COL[11001] = 1'b0;
assign COL[11002] = 1'b0;
assign COL[11003] = 1'b0;
assign COL[11004] = 1'b0;
assign COL[11005] = 1'b0;
assign COL[11006] = 1'b0;
assign COL[11007] = 1'b0;
assign COL[11008] = 1'b0;
assign COL[11009] = 1'b0;
assign COL[11010] = 1'b0;
assign COL[11011] = 1'b0;
assign COL[11012] = 1'b0;
assign COL[11013] = 1'b0;
assign COL[11014] = 1'b0;
assign COL[11015] = 1'b0;
assign COL[11016] = 1'b0;
assign COL[11017] = 1'b0;
assign COL[11018] = 1'b0;
assign COL[11019] = 1'b0;
assign COL[11020] = 1'b0;
assign COL[11021] = 1'b0;
assign COL[11022] = 1'b0;
assign COL[11023] = 1'b0;
assign COL[11024] = 1'b0;
assign COL[11025] = 1'b0;
assign COL[11026] = 1'b0;
assign COL[11027] = 1'b0;
assign COL[11028] = 1'b0;
assign COL[11029] = 1'b0;
assign COL[11030] = 1'b0;
assign COL[11031] = 1'b0;
assign COL[11032] = 1'b0;
assign COL[11033] = 1'b0;
assign COL[11034] = 1'b0;
assign COL[11035] = 1'b0;
assign COL[11036] = 1'b0;
assign COL[11037] = 1'b0;
assign COL[11038] = 1'b0;
assign COL[11039] = 1'b0;
assign COL[11040] = 1'b0;
assign COL[11041] = 1'b1;
assign COL[11042] = 1'b1;
assign COL[11043] = 1'b1;
assign COL[11044] = 1'b1;
assign COL[11045] = 1'b0;
assign COL[11046] = 1'b0;
assign COL[11047] = 1'b0;
assign COL[11048] = 1'b0;
assign COL[11049] = 1'b0;
assign COL[11050] = 1'b0;
assign COL[11051] = 1'b0;
assign COL[11052] = 1'b0;
assign COL[11053] = 1'b0;
assign COL[11054] = 1'b0;
assign COL[11055] = 1'b0;
assign COL[11056] = 1'b0;
assign COL[11057] = 1'b0;
assign COL[11058] = 1'b0;
assign COL[11059] = 1'b0;
assign COL[11060] = 1'b0;
assign COL[11061] = 1'b0;
assign COL[11062] = 1'b0;
assign COL[11063] = 1'b0;
assign COL[11064] = 1'b0;
assign COL[11065] = 1'b0;
assign COL[11066] = 1'b0;
assign COL[11067] = 1'b0;
assign COL[11068] = 1'b0;
assign COL[11069] = 1'b0;
assign COL[11070] = 1'b0;
assign COL[11071] = 1'b0;
assign COL[11072] = 1'b0;
assign COL[11073] = 1'b0;
assign COL[11074] = 1'b0;
assign COL[11075] = 1'b0;
assign COL[11076] = 1'b0;
assign COL[11077] = 1'b0;
assign COL[11078] = 1'b0;
assign COL[11079] = 1'b0;
assign COL[11080] = 1'b0;
assign COL[11081] = 1'b0;
assign COL[11082] = 1'b0;
assign COL[11083] = 1'b0;
assign COL[11084] = 1'b0;
assign COL[11085] = 1'b1;
assign COL[11086] = 1'b1;
assign COL[11087] = 1'b1;
assign COL[11088] = 1'b1;
assign COL[11089] = 1'b0;
assign COL[11090] = 1'b0;
assign COL[11091] = 1'b0;
assign COL[11092] = 1'b0;
assign COL[11093] = 1'b0;
assign COL[11094] = 1'b0;
assign COL[11095] = 1'b0;
assign COL[11096] = 1'b0;
assign COL[11097] = 1'b0;
assign COL[11098] = 1'b0;
assign COL[11099] = 1'b0;
assign COL[11100] = 1'b0;
assign COL[11101] = 1'b0;
assign COL[11102] = 1'b0;
assign COL[11103] = 1'b0;
assign COL[11104] = 1'b0;
assign COL[11105] = 1'b0;
assign COL[11106] = 1'b0;
assign COL[11107] = 1'b0;
assign COL[11108] = 1'b0;
assign COL[11109] = 1'b0;
assign COL[11110] = 1'b0;
assign COL[11111] = 1'b0;
assign COL[11112] = 1'b0;
assign COL[11113] = 1'b0;
assign COL[11114] = 1'b0;
assign COL[11115] = 1'b0;
assign COL[11116] = 1'b0;
assign COL[11117] = 1'b0;
assign COL[11118] = 1'b0;
assign COL[11119] = 1'b0;
assign COL[11120] = 1'b0;
assign COL[11121] = 1'b0;
assign COL[11122] = 1'b0;
assign COL[11123] = 1'b0;
assign COL[11124] = 1'b0;
assign COL[11125] = 1'b0;
assign COL[11126] = 1'b0;
assign COL[11127] = 1'b0;
assign COL[11128] = 1'b0;
assign COL[11129] = 1'b0;
assign COL[11130] = 1'b1;
assign COL[11131] = 1'b1;
assign COL[11132] = 1'b1;
assign COL[11133] = 1'b1;
assign COL[11134] = 1'b1;
assign COL[11135] = 1'b0;
assign COL[11136] = 1'b0;
assign COL[11137] = 1'b0;
assign COL[11138] = 1'b0;
assign COL[11139] = 1'b0;
assign COL[11140] = 1'b0;
assign COL[11141] = 1'b0;
assign COL[11142] = 1'b0;
assign COL[11143] = 1'b0;
assign COL[11144] = 1'b0;
assign COL[11145] = 1'b0;
assign COL[11146] = 1'b0;
assign COL[11147] = 1'b0;
assign COL[11148] = 1'b0;
assign COL[11149] = 1'b0;
assign COL[11150] = 1'b0;
assign COL[11151] = 1'b0;
assign COL[11152] = 1'b0;
assign COL[11153] = 1'b0;
assign COL[11154] = 1'b0;
assign COL[11155] = 1'b0;
assign COL[11156] = 1'b0;
assign COL[11157] = 1'b0;
assign COL[11158] = 1'b0;
assign COL[11159] = 1'b0;
assign COL[11160] = 1'b0;
assign COL[11161] = 1'b0;
assign COL[11162] = 1'b0;
assign COL[11163] = 1'b0;
assign COL[11164] = 1'b0;
assign COL[11165] = 1'b0;
assign COL[11166] = 1'b0;
assign COL[11167] = 1'b0;
assign COL[11168] = 1'b0;
assign COL[11169] = 1'b0;
assign COL[11170] = 1'b0;
assign COL[11171] = 1'b0;
assign COL[11172] = 1'b0;
assign COL[11173] = 1'b0;
assign COL[11174] = 1'b0;
assign COL[11175] = 1'b0;
assign COL[11176] = 1'b0;
assign COL[11177] = 1'b0;
assign COL[11178] = 1'b0;
assign COL[11179] = 1'b0;
assign COL[11180] = 1'b0;
assign COL[11181] = 1'b0;
assign COL[11182] = 1'b0;
assign COL[11183] = 1'b0;
assign COL[11184] = 1'b0;
assign COL[11185] = 1'b0;
assign COL[11186] = 1'b0;
assign COL[11187] = 1'b0;
assign COL[11188] = 1'b0;
assign COL[11189] = 1'b0;
assign COL[11190] = 1'b0;
assign COL[11191] = 1'b0;
assign COL[11192] = 1'b0;
assign COL[11193] = 1'b0;
assign COL[11194] = 1'b0;
assign COL[11195] = 1'b0;
assign COL[11196] = 1'b0;
assign COL[11197] = 1'b0;
assign COL[11198] = 1'b0;
assign COL[11199] = 1'b0;
assign COL[11200] = 1'b0;
assign COL[11201] = 1'b1;
assign COL[11202] = 1'b1;
assign COL[11203] = 1'b1;
assign COL[11204] = 1'b1;
assign COL[11205] = 1'b0;
assign COL[11206] = 1'b0;
assign COL[11207] = 1'b0;
assign COL[11208] = 1'b0;
assign COL[11209] = 1'b0;
assign COL[11210] = 1'b0;
assign COL[11211] = 1'b0;
assign COL[11212] = 1'b0;
assign COL[11213] = 1'b0;
assign COL[11214] = 1'b0;
assign COL[11215] = 1'b0;
assign COL[11216] = 1'b0;
assign COL[11217] = 1'b0;
assign COL[11218] = 1'b0;
assign COL[11219] = 1'b0;
assign COL[11220] = 1'b0;
assign COL[11221] = 1'b0;
assign COL[11222] = 1'b0;
assign COL[11223] = 1'b0;
assign COL[11224] = 1'b0;
assign COL[11225] = 1'b0;
assign COL[11226] = 1'b0;
assign COL[11227] = 1'b0;
assign COL[11228] = 1'b0;
assign COL[11229] = 1'b0;
assign COL[11230] = 1'b0;
assign COL[11231] = 1'b0;
assign COL[11232] = 1'b0;
assign COL[11233] = 1'b0;
assign COL[11234] = 1'b0;
assign COL[11235] = 1'b0;
assign COL[11236] = 1'b0;
assign COL[11237] = 1'b0;
assign COL[11238] = 1'b0;
assign COL[11239] = 1'b0;
assign COL[11240] = 1'b0;
assign COL[11241] = 1'b0;
assign COL[11242] = 1'b0;
assign COL[11243] = 1'b0;
assign COL[11244] = 1'b0;
assign COL[11245] = 1'b1;
assign COL[11246] = 1'b1;
assign COL[11247] = 1'b1;
assign COL[11248] = 1'b1;
assign COL[11249] = 1'b0;
assign COL[11250] = 1'b0;
assign COL[11251] = 1'b0;
assign COL[11252] = 1'b0;
assign COL[11253] = 1'b0;
assign COL[11254] = 1'b0;
assign COL[11255] = 1'b0;
assign COL[11256] = 1'b0;
assign COL[11257] = 1'b0;
assign COL[11258] = 1'b0;
assign COL[11259] = 1'b0;
assign COL[11260] = 1'b0;
assign COL[11261] = 1'b0;
assign COL[11262] = 1'b0;
assign COL[11263] = 1'b0;
assign COL[11264] = 1'b0;
assign COL[11265] = 1'b0;
assign COL[11266] = 1'b0;
assign COL[11267] = 1'b0;
assign COL[11268] = 1'b0;
assign COL[11269] = 1'b0;
assign COL[11270] = 1'b0;
assign COL[11271] = 1'b0;
assign COL[11272] = 1'b0;
assign COL[11273] = 1'b0;
assign COL[11274] = 1'b0;
assign COL[11275] = 1'b0;
assign COL[11276] = 1'b0;
assign COL[11277] = 1'b0;
assign COL[11278] = 1'b0;
assign COL[11279] = 1'b0;
assign COL[11280] = 1'b0;
assign COL[11281] = 1'b0;
assign COL[11282] = 1'b0;
assign COL[11283] = 1'b0;
assign COL[11284] = 1'b0;
assign COL[11285] = 1'b0;
assign COL[11286] = 1'b0;
assign COL[11287] = 1'b0;
assign COL[11288] = 1'b0;
assign COL[11289] = 1'b0;
assign COL[11290] = 1'b1;
assign COL[11291] = 1'b1;
assign COL[11292] = 1'b1;
assign COL[11293] = 1'b1;
assign COL[11294] = 1'b1;
assign COL[11295] = 1'b0;
assign COL[11296] = 1'b0;
assign COL[11297] = 1'b0;
assign COL[11298] = 1'b0;
assign COL[11299] = 1'b0;
assign COL[11300] = 1'b0;
assign COL[11301] = 1'b0;
assign COL[11302] = 1'b0;
assign COL[11303] = 1'b0;
assign COL[11304] = 1'b0;
assign COL[11305] = 1'b0;
assign COL[11306] = 1'b0;
assign COL[11307] = 1'b0;
assign COL[11308] = 1'b0;
assign COL[11309] = 1'b0;
assign COL[11310] = 1'b0;
assign COL[11311] = 1'b0;
assign COL[11312] = 1'b0;
assign COL[11313] = 1'b0;
assign COL[11314] = 1'b0;
assign COL[11315] = 1'b0;
assign COL[11316] = 1'b0;
assign COL[11317] = 1'b0;
assign COL[11318] = 1'b0;
assign COL[11319] = 1'b0;
assign COL[11320] = 1'b0;
assign COL[11321] = 1'b0;
assign COL[11322] = 1'b0;
assign COL[11323] = 1'b0;
assign COL[11324] = 1'b0;
assign COL[11325] = 1'b0;
assign COL[11326] = 1'b0;
assign COL[11327] = 1'b0;
assign COL[11328] = 1'b0;
assign COL[11329] = 1'b0;
assign COL[11330] = 1'b0;
assign COL[11331] = 1'b0;
assign COL[11332] = 1'b0;
assign COL[11333] = 1'b0;
assign COL[11334] = 1'b0;
assign COL[11335] = 1'b0;
assign COL[11336] = 1'b0;
assign COL[11337] = 1'b0;
assign COL[11338] = 1'b0;
assign COL[11339] = 1'b0;
assign COL[11340] = 1'b0;
assign COL[11341] = 1'b0;
assign COL[11342] = 1'b0;
assign COL[11343] = 1'b0;
assign COL[11344] = 1'b0;
assign COL[11345] = 1'b0;
assign COL[11346] = 1'b0;
assign COL[11347] = 1'b0;
assign COL[11348] = 1'b0;
assign COL[11349] = 1'b0;
assign COL[11350] = 1'b0;
assign COL[11351] = 1'b0;
assign COL[11352] = 1'b0;
assign COL[11353] = 1'b0;
assign COL[11354] = 1'b0;
assign COL[11355] = 1'b0;
assign COL[11356] = 1'b0;
assign COL[11357] = 1'b0;
assign COL[11358] = 1'b0;
assign COL[11359] = 1'b0;
assign COL[11360] = 1'b0;
assign COL[11361] = 1'b1;
assign COL[11362] = 1'b1;
assign COL[11363] = 1'b1;
assign COL[11364] = 1'b1;
assign COL[11365] = 1'b0;
assign COL[11366] = 1'b0;
assign COL[11367] = 1'b0;
assign COL[11368] = 1'b0;
assign COL[11369] = 1'b0;
assign COL[11370] = 1'b0;
assign COL[11371] = 1'b0;
assign COL[11372] = 1'b0;
assign COL[11373] = 1'b0;
assign COL[11374] = 1'b0;
assign COL[11375] = 1'b0;
assign COL[11376] = 1'b0;
assign COL[11377] = 1'b0;
assign COL[11378] = 1'b0;
assign COL[11379] = 1'b0;
assign COL[11380] = 1'b0;
assign COL[11381] = 1'b0;
assign COL[11382] = 1'b0;
assign COL[11383] = 1'b0;
assign COL[11384] = 1'b0;
assign COL[11385] = 1'b0;
assign COL[11386] = 1'b0;
assign COL[11387] = 1'b0;
assign COL[11388] = 1'b0;
assign COL[11389] = 1'b0;
assign COL[11390] = 1'b0;
assign COL[11391] = 1'b0;
assign COL[11392] = 1'b0;
assign COL[11393] = 1'b0;
assign COL[11394] = 1'b0;
assign COL[11395] = 1'b0;
assign COL[11396] = 1'b0;
assign COL[11397] = 1'b0;
assign COL[11398] = 1'b0;
assign COL[11399] = 1'b0;
assign COL[11400] = 1'b0;
assign COL[11401] = 1'b0;
assign COL[11402] = 1'b0;
assign COL[11403] = 1'b0;
assign COL[11404] = 1'b0;
assign COL[11405] = 1'b1;
assign COL[11406] = 1'b1;
assign COL[11407] = 1'b1;
assign COL[11408] = 1'b1;
assign COL[11409] = 1'b0;
assign COL[11410] = 1'b0;
assign COL[11411] = 1'b0;
assign COL[11412] = 1'b0;
assign COL[11413] = 1'b0;
assign COL[11414] = 1'b0;
assign COL[11415] = 1'b0;
assign COL[11416] = 1'b0;
assign COL[11417] = 1'b0;
assign COL[11418] = 1'b0;
assign COL[11419] = 1'b0;
assign COL[11420] = 1'b0;
assign COL[11421] = 1'b0;
assign COL[11422] = 1'b0;
assign COL[11423] = 1'b0;
assign COL[11424] = 1'b0;
assign COL[11425] = 1'b0;
assign COL[11426] = 1'b0;
assign COL[11427] = 1'b0;
assign COL[11428] = 1'b0;
assign COL[11429] = 1'b0;
assign COL[11430] = 1'b0;
assign COL[11431] = 1'b0;
assign COL[11432] = 1'b0;
assign COL[11433] = 1'b0;
assign COL[11434] = 1'b0;
assign COL[11435] = 1'b0;
assign COL[11436] = 1'b0;
assign COL[11437] = 1'b0;
assign COL[11438] = 1'b0;
assign COL[11439] = 1'b0;
assign COL[11440] = 1'b0;
assign COL[11441] = 1'b0;
assign COL[11442] = 1'b0;
assign COL[11443] = 1'b0;
assign COL[11444] = 1'b0;
assign COL[11445] = 1'b0;
assign COL[11446] = 1'b0;
assign COL[11447] = 1'b0;
assign COL[11448] = 1'b0;
assign COL[11449] = 1'b0;
assign COL[11450] = 1'b1;
assign COL[11451] = 1'b1;
assign COL[11452] = 1'b1;
assign COL[11453] = 1'b1;
assign COL[11454] = 1'b1;
assign COL[11455] = 1'b0;
assign COL[11456] = 1'b0;
assign COL[11457] = 1'b0;
assign COL[11458] = 1'b0;
assign COL[11459] = 1'b0;
assign COL[11460] = 1'b0;
assign COL[11461] = 1'b0;
assign COL[11462] = 1'b0;
assign COL[11463] = 1'b0;
assign COL[11464] = 1'b0;
assign COL[11465] = 1'b0;
assign COL[11466] = 1'b0;
assign COL[11467] = 1'b0;
assign COL[11468] = 1'b0;
assign COL[11469] = 1'b0;
assign COL[11470] = 1'b0;
assign COL[11471] = 1'b0;
assign COL[11472] = 1'b0;
assign COL[11473] = 1'b0;
assign COL[11474] = 1'b0;
assign COL[11475] = 1'b0;
assign COL[11476] = 1'b0;
assign COL[11477] = 1'b0;
assign COL[11478] = 1'b0;
assign COL[11479] = 1'b0;
assign COL[11480] = 1'b0;
assign COL[11481] = 1'b0;
assign COL[11482] = 1'b0;
assign COL[11483] = 1'b0;
assign COL[11484] = 1'b0;
assign COL[11485] = 1'b0;
assign COL[11486] = 1'b0;
assign COL[11487] = 1'b0;
assign COL[11488] = 1'b0;
assign COL[11489] = 1'b0;
assign COL[11490] = 1'b0;
assign COL[11491] = 1'b0;
assign COL[11492] = 1'b0;
assign COL[11493] = 1'b0;
assign COL[11494] = 1'b0;
assign COL[11495] = 1'b0;
assign COL[11496] = 1'b0;
assign COL[11497] = 1'b0;
assign COL[11498] = 1'b0;
assign COL[11499] = 1'b0;
assign COL[11500] = 1'b0;
assign COL[11501] = 1'b0;
assign COL[11502] = 1'b0;
assign COL[11503] = 1'b0;
assign COL[11504] = 1'b0;
assign COL[11505] = 1'b0;
assign COL[11506] = 1'b0;
assign COL[11507] = 1'b0;
assign COL[11508] = 1'b0;
assign COL[11509] = 1'b0;
assign COL[11510] = 1'b0;
assign COL[11511] = 1'b0;
assign COL[11512] = 1'b0;
assign COL[11513] = 1'b0;
assign COL[11514] = 1'b0;
assign COL[11515] = 1'b0;
assign COL[11516] = 1'b0;
assign COL[11517] = 1'b0;
assign COL[11518] = 1'b0;
assign COL[11519] = 1'b0;
assign COL[11520] = 1'b0;
assign COL[11521] = 1'b1;
assign COL[11522] = 1'b1;
assign COL[11523] = 1'b1;
assign COL[11524] = 1'b1;
assign COL[11525] = 1'b0;
assign COL[11526] = 1'b0;
assign COL[11527] = 1'b0;
assign COL[11528] = 1'b0;
assign COL[11529] = 1'b0;
assign COL[11530] = 1'b0;
assign COL[11531] = 1'b0;
assign COL[11532] = 1'b0;
assign COL[11533] = 1'b0;
assign COL[11534] = 1'b0;
assign COL[11535] = 1'b0;
assign COL[11536] = 1'b0;
assign COL[11537] = 1'b0;
assign COL[11538] = 1'b0;
assign COL[11539] = 1'b0;
assign COL[11540] = 1'b0;
assign COL[11541] = 1'b0;
assign COL[11542] = 1'b0;
assign COL[11543] = 1'b0;
assign COL[11544] = 1'b0;
assign COL[11545] = 1'b0;
assign COL[11546] = 1'b0;
assign COL[11547] = 1'b0;
assign COL[11548] = 1'b0;
assign COL[11549] = 1'b0;
assign COL[11550] = 1'b0;
assign COL[11551] = 1'b0;
assign COL[11552] = 1'b0;
assign COL[11553] = 1'b0;
assign COL[11554] = 1'b0;
assign COL[11555] = 1'b0;
assign COL[11556] = 1'b0;
assign COL[11557] = 1'b0;
assign COL[11558] = 1'b0;
assign COL[11559] = 1'b0;
assign COL[11560] = 1'b0;
assign COL[11561] = 1'b0;
assign COL[11562] = 1'b0;
assign COL[11563] = 1'b0;
assign COL[11564] = 1'b0;
assign COL[11565] = 1'b1;
assign COL[11566] = 1'b1;
assign COL[11567] = 1'b1;
assign COL[11568] = 1'b1;
assign COL[11569] = 1'b0;
assign COL[11570] = 1'b0;
assign COL[11571] = 1'b0;
assign COL[11572] = 1'b0;
assign COL[11573] = 1'b0;
assign COL[11574] = 1'b0;
assign COL[11575] = 1'b0;
assign COL[11576] = 1'b0;
assign COL[11577] = 1'b0;
assign COL[11578] = 1'b0;
assign COL[11579] = 1'b0;
assign COL[11580] = 1'b0;
assign COL[11581] = 1'b0;
assign COL[11582] = 1'b0;
assign COL[11583] = 1'b0;
assign COL[11584] = 1'b0;
assign COL[11585] = 1'b0;
assign COL[11586] = 1'b0;
assign COL[11587] = 1'b0;
assign COL[11588] = 1'b0;
assign COL[11589] = 1'b0;
assign COL[11590] = 1'b0;
assign COL[11591] = 1'b0;
assign COL[11592] = 1'b0;
assign COL[11593] = 1'b0;
assign COL[11594] = 1'b0;
assign COL[11595] = 1'b0;
assign COL[11596] = 1'b0;
assign COL[11597] = 1'b0;
assign COL[11598] = 1'b0;
assign COL[11599] = 1'b0;
assign COL[11600] = 1'b0;
assign COL[11601] = 1'b0;
assign COL[11602] = 1'b0;
assign COL[11603] = 1'b0;
assign COL[11604] = 1'b0;
assign COL[11605] = 1'b0;
assign COL[11606] = 1'b0;
assign COL[11607] = 1'b0;
assign COL[11608] = 1'b0;
assign COL[11609] = 1'b0;
assign COL[11610] = 1'b1;
assign COL[11611] = 1'b1;
assign COL[11612] = 1'b1;
assign COL[11613] = 1'b1;
assign COL[11614] = 1'b1;
assign COL[11615] = 1'b0;
assign COL[11616] = 1'b0;
assign COL[11617] = 1'b0;
assign COL[11618] = 1'b0;
assign COL[11619] = 1'b0;
assign COL[11620] = 1'b0;
assign COL[11621] = 1'b0;
assign COL[11622] = 1'b0;
assign COL[11623] = 1'b0;
assign COL[11624] = 1'b0;
assign COL[11625] = 1'b0;
assign COL[11626] = 1'b0;
assign COL[11627] = 1'b0;
assign COL[11628] = 1'b0;
assign COL[11629] = 1'b0;
assign COL[11630] = 1'b0;
assign COL[11631] = 1'b0;
assign COL[11632] = 1'b0;
assign COL[11633] = 1'b0;
assign COL[11634] = 1'b0;
assign COL[11635] = 1'b0;
assign COL[11636] = 1'b0;
assign COL[11637] = 1'b0;
assign COL[11638] = 1'b0;
assign COL[11639] = 1'b0;
assign COL[11640] = 1'b0;
assign COL[11641] = 1'b0;
assign COL[11642] = 1'b0;
assign COL[11643] = 1'b0;
assign COL[11644] = 1'b0;
assign COL[11645] = 1'b0;
assign COL[11646] = 1'b0;
assign COL[11647] = 1'b0;
assign COL[11648] = 1'b0;
assign COL[11649] = 1'b0;
assign COL[11650] = 1'b0;
assign COL[11651] = 1'b0;
assign COL[11652] = 1'b0;
assign COL[11653] = 1'b0;
assign COL[11654] = 1'b0;
assign COL[11655] = 1'b0;
assign COL[11656] = 1'b0;
assign COL[11657] = 1'b0;
assign COL[11658] = 1'b0;
assign COL[11659] = 1'b0;
assign COL[11660] = 1'b0;
assign COL[11661] = 1'b0;
assign COL[11662] = 1'b0;
assign COL[11663] = 1'b0;
assign COL[11664] = 1'b0;
assign COL[11665] = 1'b0;
assign COL[11666] = 1'b0;
assign COL[11667] = 1'b0;
assign COL[11668] = 1'b0;
assign COL[11669] = 1'b0;
assign COL[11670] = 1'b0;
assign COL[11671] = 1'b0;
assign COL[11672] = 1'b0;
assign COL[11673] = 1'b0;
assign COL[11674] = 1'b0;
assign COL[11675] = 1'b0;
assign COL[11676] = 1'b0;
assign COL[11677] = 1'b0;
assign COL[11678] = 1'b0;
assign COL[11679] = 1'b0;
assign COL[11680] = 1'b0;
assign COL[11681] = 1'b1;
assign COL[11682] = 1'b1;
assign COL[11683] = 1'b1;
assign COL[11684] = 1'b1;
assign COL[11685] = 1'b0;
assign COL[11686] = 1'b0;
assign COL[11687] = 1'b0;
assign COL[11688] = 1'b0;
assign COL[11689] = 1'b0;
assign COL[11690] = 1'b0;
assign COL[11691] = 1'b0;
assign COL[11692] = 1'b0;
assign COL[11693] = 1'b0;
assign COL[11694] = 1'b0;
assign COL[11695] = 1'b0;
assign COL[11696] = 1'b0;
assign COL[11697] = 1'b0;
assign COL[11698] = 1'b0;
assign COL[11699] = 1'b0;
assign COL[11700] = 1'b0;
assign COL[11701] = 1'b0;
assign COL[11702] = 1'b0;
assign COL[11703] = 1'b0;
assign COL[11704] = 1'b0;
assign COL[11705] = 1'b0;
assign COL[11706] = 1'b0;
assign COL[11707] = 1'b0;
assign COL[11708] = 1'b0;
assign COL[11709] = 1'b0;
assign COL[11710] = 1'b0;
assign COL[11711] = 1'b0;
assign COL[11712] = 1'b0;
assign COL[11713] = 1'b0;
assign COL[11714] = 1'b0;
assign COL[11715] = 1'b0;
assign COL[11716] = 1'b0;
assign COL[11717] = 1'b0;
assign COL[11718] = 1'b0;
assign COL[11719] = 1'b0;
assign COL[11720] = 1'b0;
assign COL[11721] = 1'b0;
assign COL[11722] = 1'b0;
assign COL[11723] = 1'b0;
assign COL[11724] = 1'b0;
assign COL[11725] = 1'b1;
assign COL[11726] = 1'b1;
assign COL[11727] = 1'b1;
assign COL[11728] = 1'b1;
assign COL[11729] = 1'b0;
assign COL[11730] = 1'b0;
assign COL[11731] = 1'b0;
assign COL[11732] = 1'b0;
assign COL[11733] = 1'b0;
assign COL[11734] = 1'b0;
assign COL[11735] = 1'b0;
assign COL[11736] = 1'b0;
assign COL[11737] = 1'b0;
assign COL[11738] = 1'b0;
assign COL[11739] = 1'b0;
assign COL[11740] = 1'b0;
assign COL[11741] = 1'b0;
assign COL[11742] = 1'b0;
assign COL[11743] = 1'b0;
assign COL[11744] = 1'b0;
assign COL[11745] = 1'b0;
assign COL[11746] = 1'b0;
assign COL[11747] = 1'b0;
assign COL[11748] = 1'b0;
assign COL[11749] = 1'b0;
assign COL[11750] = 1'b0;
assign COL[11751] = 1'b0;
assign COL[11752] = 1'b0;
assign COL[11753] = 1'b0;
assign COL[11754] = 1'b0;
assign COL[11755] = 1'b0;
assign COL[11756] = 1'b0;
assign COL[11757] = 1'b0;
assign COL[11758] = 1'b0;
assign COL[11759] = 1'b0;
assign COL[11760] = 1'b0;
assign COL[11761] = 1'b0;
assign COL[11762] = 1'b0;
assign COL[11763] = 1'b0;
assign COL[11764] = 1'b0;
assign COL[11765] = 1'b0;
assign COL[11766] = 1'b0;
assign COL[11767] = 1'b0;
assign COL[11768] = 1'b0;
assign COL[11769] = 1'b0;
assign COL[11770] = 1'b1;
assign COL[11771] = 1'b1;
assign COL[11772] = 1'b1;
assign COL[11773] = 1'b1;
assign COL[11774] = 1'b1;
assign COL[11775] = 1'b0;
assign COL[11776] = 1'b0;
assign COL[11777] = 1'b0;
assign COL[11778] = 1'b0;
assign COL[11779] = 1'b0;
assign COL[11780] = 1'b0;
assign COL[11781] = 1'b0;
assign COL[11782] = 1'b0;
assign COL[11783] = 1'b0;
assign COL[11784] = 1'b0;
assign COL[11785] = 1'b0;
assign COL[11786] = 1'b0;
assign COL[11787] = 1'b0;
assign COL[11788] = 1'b0;
assign COL[11789] = 1'b0;
assign COL[11790] = 1'b0;
assign COL[11791] = 1'b0;
assign COL[11792] = 1'b0;
assign COL[11793] = 1'b0;
assign COL[11794] = 1'b0;
assign COL[11795] = 1'b0;
assign COL[11796] = 1'b0;
assign COL[11797] = 1'b0;
assign COL[11798] = 1'b0;
assign COL[11799] = 1'b0;
assign COL[11800] = 1'b0;
assign COL[11801] = 1'b0;
assign COL[11802] = 1'b0;
assign COL[11803] = 1'b0;
assign COL[11804] = 1'b0;
assign COL[11805] = 1'b0;
assign COL[11806] = 1'b0;
assign COL[11807] = 1'b0;
assign COL[11808] = 1'b0;
assign COL[11809] = 1'b0;
assign COL[11810] = 1'b0;
assign COL[11811] = 1'b0;
assign COL[11812] = 1'b0;
assign COL[11813] = 1'b0;
assign COL[11814] = 1'b0;
assign COL[11815] = 1'b0;
assign COL[11816] = 1'b0;
assign COL[11817] = 1'b0;
assign COL[11818] = 1'b0;
assign COL[11819] = 1'b0;
assign COL[11820] = 1'b0;
assign COL[11821] = 1'b0;
assign COL[11822] = 1'b0;
assign COL[11823] = 1'b0;
assign COL[11824] = 1'b0;
assign COL[11825] = 1'b0;
assign COL[11826] = 1'b0;
assign COL[11827] = 1'b0;
assign COL[11828] = 1'b0;
assign COL[11829] = 1'b0;
assign COL[11830] = 1'b0;
assign COL[11831] = 1'b0;
assign COL[11832] = 1'b0;
assign COL[11833] = 1'b0;
assign COL[11834] = 1'b0;
assign COL[11835] = 1'b0;
assign COL[11836] = 1'b0;
assign COL[11837] = 1'b0;
assign COL[11838] = 1'b0;
assign COL[11839] = 1'b0;
assign COL[11840] = 1'b0;
assign COL[11841] = 1'b1;
assign COL[11842] = 1'b1;
assign COL[11843] = 1'b1;
assign COL[11844] = 1'b1;
assign COL[11845] = 1'b0;
assign COL[11846] = 1'b0;
assign COL[11847] = 1'b0;
assign COL[11848] = 1'b0;
assign COL[11849] = 1'b0;
assign COL[11850] = 1'b0;
assign COL[11851] = 1'b0;
assign COL[11852] = 1'b0;
assign COL[11853] = 1'b0;
assign COL[11854] = 1'b0;
assign COL[11855] = 1'b0;
assign COL[11856] = 1'b0;
assign COL[11857] = 1'b0;
assign COL[11858] = 1'b0;
assign COL[11859] = 1'b0;
assign COL[11860] = 1'b0;
assign COL[11861] = 1'b0;
assign COL[11862] = 1'b0;
assign COL[11863] = 1'b0;
assign COL[11864] = 1'b0;
assign COL[11865] = 1'b0;
assign COL[11866] = 1'b0;
assign COL[11867] = 1'b0;
assign COL[11868] = 1'b0;
assign COL[11869] = 1'b0;
assign COL[11870] = 1'b0;
assign COL[11871] = 1'b0;
assign COL[11872] = 1'b0;
assign COL[11873] = 1'b0;
assign COL[11874] = 1'b0;
assign COL[11875] = 1'b0;
assign COL[11876] = 1'b0;
assign COL[11877] = 1'b0;
assign COL[11878] = 1'b0;
assign COL[11879] = 1'b0;
assign COL[11880] = 1'b0;
assign COL[11881] = 1'b0;
assign COL[11882] = 1'b0;
assign COL[11883] = 1'b0;
assign COL[11884] = 1'b0;
assign COL[11885] = 1'b1;
assign COL[11886] = 1'b1;
assign COL[11887] = 1'b1;
assign COL[11888] = 1'b1;
assign COL[11889] = 1'b0;
assign COL[11890] = 1'b0;
assign COL[11891] = 1'b0;
assign COL[11892] = 1'b0;
assign COL[11893] = 1'b0;
assign COL[11894] = 1'b0;
assign COL[11895] = 1'b0;
assign COL[11896] = 1'b0;
assign COL[11897] = 1'b0;
assign COL[11898] = 1'b0;
assign COL[11899] = 1'b0;
assign COL[11900] = 1'b0;
assign COL[11901] = 1'b0;
assign COL[11902] = 1'b0;
assign COL[11903] = 1'b0;
assign COL[11904] = 1'b0;
assign COL[11905] = 1'b0;
assign COL[11906] = 1'b0;
assign COL[11907] = 1'b0;
assign COL[11908] = 1'b0;
assign COL[11909] = 1'b0;
assign COL[11910] = 1'b0;
assign COL[11911] = 1'b0;
assign COL[11912] = 1'b0;
assign COL[11913] = 1'b0;
assign COL[11914] = 1'b0;
assign COL[11915] = 1'b0;
assign COL[11916] = 1'b0;
assign COL[11917] = 1'b0;
assign COL[11918] = 1'b0;
assign COL[11919] = 1'b0;
assign COL[11920] = 1'b0;
assign COL[11921] = 1'b0;
assign COL[11922] = 1'b0;
assign COL[11923] = 1'b0;
assign COL[11924] = 1'b0;
assign COL[11925] = 1'b0;
assign COL[11926] = 1'b0;
assign COL[11927] = 1'b0;
assign COL[11928] = 1'b0;
assign COL[11929] = 1'b0;
assign COL[11930] = 1'b1;
assign COL[11931] = 1'b1;
assign COL[11932] = 1'b1;
assign COL[11933] = 1'b1;
assign COL[11934] = 1'b1;
assign COL[11935] = 1'b0;
assign COL[11936] = 1'b0;
assign COL[11937] = 1'b0;
assign COL[11938] = 1'b0;
assign COL[11939] = 1'b0;
assign COL[11940] = 1'b0;
assign COL[11941] = 1'b0;
assign COL[11942] = 1'b0;
assign COL[11943] = 1'b0;
assign COL[11944] = 1'b0;
assign COL[11945] = 1'b0;
assign COL[11946] = 1'b0;
assign COL[11947] = 1'b0;
assign COL[11948] = 1'b0;
assign COL[11949] = 1'b0;
assign COL[11950] = 1'b0;
assign COL[11951] = 1'b0;
assign COL[11952] = 1'b0;
assign COL[11953] = 1'b0;
assign COL[11954] = 1'b0;
assign COL[11955] = 1'b0;
assign COL[11956] = 1'b0;
assign COL[11957] = 1'b0;
assign COL[11958] = 1'b0;
assign COL[11959] = 1'b0;
assign COL[11960] = 1'b0;
assign COL[11961] = 1'b0;
assign COL[11962] = 1'b0;
assign COL[11963] = 1'b0;
assign COL[11964] = 1'b0;
assign COL[11965] = 1'b0;
assign COL[11966] = 1'b0;
assign COL[11967] = 1'b0;
assign COL[11968] = 1'b0;
assign COL[11969] = 1'b0;
assign COL[11970] = 1'b0;
assign COL[11971] = 1'b0;
assign COL[11972] = 1'b0;
assign COL[11973] = 1'b0;
assign COL[11974] = 1'b0;
assign COL[11975] = 1'b0;
assign COL[11976] = 1'b0;
assign COL[11977] = 1'b0;
assign COL[11978] = 1'b0;
assign COL[11979] = 1'b0;
assign COL[11980] = 1'b0;
assign COL[11981] = 1'b0;
assign COL[11982] = 1'b0;
assign COL[11983] = 1'b0;
assign COL[11984] = 1'b0;
assign COL[11985] = 1'b0;
assign COL[11986] = 1'b0;
assign COL[11987] = 1'b0;
assign COL[11988] = 1'b0;
assign COL[11989] = 1'b0;
assign COL[11990] = 1'b0;
assign COL[11991] = 1'b0;
assign COL[11992] = 1'b0;
assign COL[11993] = 1'b0;
assign COL[11994] = 1'b0;
assign COL[11995] = 1'b0;
assign COL[11996] = 1'b0;
assign COL[11997] = 1'b0;
assign COL[11998] = 1'b0;
assign COL[11999] = 1'b0;
assign COL[12000] = 1'b0;
assign COL[12001] = 1'b1;
assign COL[12002] = 1'b1;
assign COL[12003] = 1'b1;
assign COL[12004] = 1'b1;
assign COL[12005] = 1'b0;
assign COL[12006] = 1'b0;
assign COL[12007] = 1'b0;
assign COL[12008] = 1'b0;
assign COL[12009] = 1'b0;
assign COL[12010] = 1'b0;
assign COL[12011] = 1'b0;
assign COL[12012] = 1'b0;
assign COL[12013] = 1'b0;
assign COL[12014] = 1'b0;
assign COL[12015] = 1'b0;
assign COL[12016] = 1'b0;
assign COL[12017] = 1'b0;
assign COL[12018] = 1'b0;
assign COL[12019] = 1'b0;
assign COL[12020] = 1'b0;
assign COL[12021] = 1'b0;
assign COL[12022] = 1'b0;
assign COL[12023] = 1'b0;
assign COL[12024] = 1'b0;
assign COL[12025] = 1'b0;
assign COL[12026] = 1'b0;
assign COL[12027] = 1'b0;
assign COL[12028] = 1'b0;
assign COL[12029] = 1'b0;
assign COL[12030] = 1'b0;
assign COL[12031] = 1'b0;
assign COL[12032] = 1'b0;
assign COL[12033] = 1'b0;
assign COL[12034] = 1'b0;
assign COL[12035] = 1'b0;
assign COL[12036] = 1'b0;
assign COL[12037] = 1'b0;
assign COL[12038] = 1'b0;
assign COL[12039] = 1'b0;
assign COL[12040] = 1'b0;
assign COL[12041] = 1'b0;
assign COL[12042] = 1'b0;
assign COL[12043] = 1'b0;
assign COL[12044] = 1'b0;
assign COL[12045] = 1'b1;
assign COL[12046] = 1'b1;
assign COL[12047] = 1'b1;
assign COL[12048] = 1'b1;
assign COL[12049] = 1'b0;
assign COL[12050] = 1'b0;
assign COL[12051] = 1'b0;
assign COL[12052] = 1'b0;
assign COL[12053] = 1'b0;
assign COL[12054] = 1'b0;
assign COL[12055] = 1'b1;
assign COL[12056] = 1'b1;
assign COL[12057] = 1'b1;
assign COL[12058] = 1'b1;
assign COL[12059] = 1'b0;
assign COL[12060] = 1'b0;
assign COL[12061] = 1'b0;
assign COL[12062] = 1'b0;
assign COL[12063] = 1'b0;
assign COL[12064] = 1'b0;
assign COL[12065] = 1'b0;
assign COL[12066] = 1'b0;
assign COL[12067] = 1'b0;
assign COL[12068] = 1'b0;
assign COL[12069] = 1'b0;
assign COL[12070] = 1'b0;
assign COL[12071] = 1'b0;
assign COL[12072] = 1'b0;
assign COL[12073] = 1'b0;
assign COL[12074] = 1'b0;
assign COL[12075] = 1'b0;
assign COL[12076] = 1'b0;
assign COL[12077] = 1'b0;
assign COL[12078] = 1'b0;
assign COL[12079] = 1'b0;
assign COL[12080] = 1'b0;
assign COL[12081] = 1'b0;
assign COL[12082] = 1'b0;
assign COL[12083] = 1'b0;
assign COL[12084] = 1'b0;
assign COL[12085] = 1'b0;
assign COL[12086] = 1'b0;
assign COL[12087] = 1'b0;
assign COL[12088] = 1'b0;
assign COL[12089] = 1'b0;
assign COL[12090] = 1'b1;
assign COL[12091] = 1'b1;
assign COL[12092] = 1'b1;
assign COL[12093] = 1'b1;
assign COL[12094] = 1'b1;
assign COL[12095] = 1'b0;
assign COL[12096] = 1'b0;
assign COL[12097] = 1'b0;
assign COL[12098] = 1'b0;
assign COL[12099] = 1'b0;
assign COL[12100] = 1'b0;
assign COL[12101] = 1'b0;
assign COL[12102] = 1'b0;
assign COL[12103] = 1'b0;
assign COL[12104] = 1'b0;
assign COL[12105] = 1'b0;
assign COL[12106] = 1'b0;
assign COL[12107] = 1'b0;
assign COL[12108] = 1'b0;
assign COL[12109] = 1'b0;
assign COL[12110] = 1'b0;
assign COL[12111] = 1'b0;
assign COL[12112] = 1'b0;
assign COL[12113] = 1'b0;
assign COL[12114] = 1'b0;
assign COL[12115] = 1'b0;
assign COL[12116] = 1'b0;
assign COL[12117] = 1'b0;
assign COL[12118] = 1'b0;
assign COL[12119] = 1'b0;
assign COL[12120] = 1'b0;
assign COL[12121] = 1'b0;
assign COL[12122] = 1'b0;
assign COL[12123] = 1'b0;
assign COL[12124] = 1'b0;
assign COL[12125] = 1'b0;
assign COL[12126] = 1'b0;
assign COL[12127] = 1'b0;
assign COL[12128] = 1'b0;
assign COL[12129] = 1'b0;
assign COL[12130] = 1'b0;
assign COL[12131] = 1'b0;
assign COL[12132] = 1'b0;
assign COL[12133] = 1'b0;
assign COL[12134] = 1'b0;
assign COL[12135] = 1'b0;
assign COL[12136] = 1'b0;
assign COL[12137] = 1'b0;
assign COL[12138] = 1'b0;
assign COL[12139] = 1'b0;
assign COL[12140] = 1'b0;
assign COL[12141] = 1'b0;
assign COL[12142] = 1'b0;
assign COL[12143] = 1'b0;
assign COL[12144] = 1'b0;
assign COL[12145] = 1'b0;
assign COL[12146] = 1'b0;
assign COL[12147] = 1'b0;
assign COL[12148] = 1'b0;
assign COL[12149] = 1'b0;
assign COL[12150] = 1'b0;
assign COL[12151] = 1'b0;
assign COL[12152] = 1'b0;
assign COL[12153] = 1'b0;
assign COL[12154] = 1'b0;
assign COL[12155] = 1'b0;
assign COL[12156] = 1'b0;
assign COL[12157] = 1'b0;
assign COL[12158] = 1'b0;
assign COL[12159] = 1'b0;
assign COL[12160] = 1'b0;
assign COL[12161] = 1'b1;
assign COL[12162] = 1'b1;
assign COL[12163] = 1'b1;
assign COL[12164] = 1'b1;
assign COL[12165] = 1'b0;
assign COL[12166] = 1'b0;
assign COL[12167] = 1'b0;
assign COL[12168] = 1'b0;
assign COL[12169] = 1'b0;
assign COL[12170] = 1'b0;
assign COL[12171] = 1'b0;
assign COL[12172] = 1'b0;
assign COL[12173] = 1'b0;
assign COL[12174] = 1'b0;
assign COL[12175] = 1'b0;
assign COL[12176] = 1'b0;
assign COL[12177] = 1'b0;
assign COL[12178] = 1'b0;
assign COL[12179] = 1'b0;
assign COL[12180] = 1'b0;
assign COL[12181] = 1'b0;
assign COL[12182] = 1'b0;
assign COL[12183] = 1'b0;
assign COL[12184] = 1'b0;
assign COL[12185] = 1'b0;
assign COL[12186] = 1'b0;
assign COL[12187] = 1'b0;
assign COL[12188] = 1'b0;
assign COL[12189] = 1'b0;
assign COL[12190] = 1'b0;
assign COL[12191] = 1'b0;
assign COL[12192] = 1'b0;
assign COL[12193] = 1'b0;
assign COL[12194] = 1'b0;
assign COL[12195] = 1'b0;
assign COL[12196] = 1'b0;
assign COL[12197] = 1'b0;
assign COL[12198] = 1'b0;
assign COL[12199] = 1'b0;
assign COL[12200] = 1'b0;
assign COL[12201] = 1'b0;
assign COL[12202] = 1'b0;
assign COL[12203] = 1'b0;
assign COL[12204] = 1'b0;
assign COL[12205] = 1'b1;
assign COL[12206] = 1'b1;
assign COL[12207] = 1'b1;
assign COL[12208] = 1'b1;
assign COL[12209] = 1'b0;
assign COL[12210] = 1'b0;
assign COL[12211] = 1'b0;
assign COL[12212] = 1'b0;
assign COL[12213] = 1'b0;
assign COL[12214] = 1'b0;
assign COL[12215] = 1'b1;
assign COL[12216] = 1'b1;
assign COL[12217] = 1'b1;
assign COL[12218] = 1'b1;
assign COL[12219] = 1'b0;
assign COL[12220] = 1'b0;
assign COL[12221] = 1'b0;
assign COL[12222] = 1'b0;
assign COL[12223] = 1'b0;
assign COL[12224] = 1'b0;
assign COL[12225] = 1'b0;
assign COL[12226] = 1'b0;
assign COL[12227] = 1'b0;
assign COL[12228] = 1'b0;
assign COL[12229] = 1'b0;
assign COL[12230] = 1'b0;
assign COL[12231] = 1'b0;
assign COL[12232] = 1'b0;
assign COL[12233] = 1'b0;
assign COL[12234] = 1'b0;
assign COL[12235] = 1'b0;
assign COL[12236] = 1'b0;
assign COL[12237] = 1'b0;
assign COL[12238] = 1'b0;
assign COL[12239] = 1'b0;
assign COL[12240] = 1'b0;
assign COL[12241] = 1'b0;
assign COL[12242] = 1'b0;
assign COL[12243] = 1'b0;
assign COL[12244] = 1'b0;
assign COL[12245] = 1'b0;
assign COL[12246] = 1'b0;
assign COL[12247] = 1'b0;
assign COL[12248] = 1'b0;
assign COL[12249] = 1'b0;
assign COL[12250] = 1'b1;
assign COL[12251] = 1'b1;
assign COL[12252] = 1'b1;
assign COL[12253] = 1'b1;
assign COL[12254] = 1'b1;
assign COL[12255] = 1'b0;
assign COL[12256] = 1'b0;
assign COL[12257] = 1'b0;
assign COL[12258] = 1'b0;
assign COL[12259] = 1'b0;
assign COL[12260] = 1'b0;
assign COL[12261] = 1'b0;
assign COL[12262] = 1'b0;
assign COL[12263] = 1'b0;
assign COL[12264] = 1'b0;
assign COL[12265] = 1'b0;
assign COL[12266] = 1'b0;
assign COL[12267] = 1'b0;
assign COL[12268] = 1'b0;
assign COL[12269] = 1'b0;
assign COL[12270] = 1'b0;
assign COL[12271] = 1'b0;
assign COL[12272] = 1'b0;
assign COL[12273] = 1'b0;
assign COL[12274] = 1'b0;
assign COL[12275] = 1'b0;
assign COL[12276] = 1'b0;
assign COL[12277] = 1'b0;
assign COL[12278] = 1'b0;
assign COL[12279] = 1'b0;
assign COL[12280] = 1'b0;
assign COL[12281] = 1'b0;
assign COL[12282] = 1'b0;
assign COL[12283] = 1'b0;
assign COL[12284] = 1'b0;
assign COL[12285] = 1'b0;
assign COL[12286] = 1'b0;
assign COL[12287] = 1'b0;
assign COL[12288] = 1'b0;
assign COL[12289] = 1'b0;
assign COL[12290] = 1'b0;
assign COL[12291] = 1'b0;
assign COL[12292] = 1'b0;
assign COL[12293] = 1'b0;
assign COL[12294] = 1'b0;
assign COL[12295] = 1'b0;
assign COL[12296] = 1'b0;
assign COL[12297] = 1'b0;
assign COL[12298] = 1'b0;
assign COL[12299] = 1'b0;
assign COL[12300] = 1'b0;
assign COL[12301] = 1'b0;
assign COL[12302] = 1'b0;
assign COL[12303] = 1'b0;
assign COL[12304] = 1'b0;
assign COL[12305] = 1'b0;
assign COL[12306] = 1'b0;
assign COL[12307] = 1'b0;
assign COL[12308] = 1'b0;
assign COL[12309] = 1'b0;
assign COL[12310] = 1'b0;
assign COL[12311] = 1'b0;
assign COL[12312] = 1'b0;
assign COL[12313] = 1'b0;
assign COL[12314] = 1'b0;
assign COL[12315] = 1'b0;
assign COL[12316] = 1'b0;
assign COL[12317] = 1'b0;
assign COL[12318] = 1'b0;
assign COL[12319] = 1'b0;
assign COL[12320] = 1'b0;
assign COL[12321] = 1'b1;
assign COL[12322] = 1'b1;
assign COL[12323] = 1'b1;
assign COL[12324] = 1'b1;
assign COL[12325] = 1'b0;
assign COL[12326] = 1'b0;
assign COL[12327] = 1'b0;
assign COL[12328] = 1'b0;
assign COL[12329] = 1'b0;
assign COL[12330] = 1'b0;
assign COL[12331] = 1'b1;
assign COL[12332] = 1'b1;
assign COL[12333] = 1'b1;
assign COL[12334] = 1'b1;
assign COL[12335] = 1'b1;
assign COL[12336] = 1'b1;
assign COL[12337] = 1'b1;
assign COL[12338] = 1'b1;
assign COL[12339] = 1'b1;
assign COL[12340] = 1'b1;
assign COL[12341] = 1'b1;
assign COL[12342] = 1'b1;
assign COL[12343] = 1'b1;
assign COL[12344] = 1'b1;
assign COL[12345] = 1'b1;
assign COL[12346] = 1'b1;
assign COL[12347] = 1'b1;
assign COL[12348] = 1'b1;
assign COL[12349] = 1'b1;
assign COL[12350] = 1'b1;
assign COL[12351] = 1'b1;
assign COL[12352] = 1'b1;
assign COL[12353] = 1'b1;
assign COL[12354] = 1'b1;
assign COL[12355] = 1'b1;
assign COL[12356] = 1'b1;
assign COL[12357] = 1'b1;
assign COL[12358] = 1'b1;
assign COL[12359] = 1'b1;
assign COL[12360] = 1'b1;
assign COL[12361] = 1'b1;
assign COL[12362] = 1'b1;
assign COL[12363] = 1'b1;
assign COL[12364] = 1'b1;
assign COL[12365] = 1'b1;
assign COL[12366] = 1'b1;
assign COL[12367] = 1'b1;
assign COL[12368] = 1'b1;
assign COL[12369] = 1'b0;
assign COL[12370] = 1'b0;
assign COL[12371] = 1'b0;
assign COL[12372] = 1'b0;
assign COL[12373] = 1'b0;
assign COL[12374] = 1'b0;
assign COL[12375] = 1'b1;
assign COL[12376] = 1'b1;
assign COL[12377] = 1'b1;
assign COL[12378] = 1'b1;
assign COL[12379] = 1'b0;
assign COL[12380] = 1'b0;
assign COL[12381] = 1'b0;
assign COL[12382] = 1'b0;
assign COL[12383] = 1'b0;
assign COL[12384] = 1'b0;
assign COL[12385] = 1'b0;
assign COL[12386] = 1'b0;
assign COL[12387] = 1'b0;
assign COL[12388] = 1'b0;
assign COL[12389] = 1'b0;
assign COL[12390] = 1'b0;
assign COL[12391] = 1'b0;
assign COL[12392] = 1'b0;
assign COL[12393] = 1'b0;
assign COL[12394] = 1'b0;
assign COL[12395] = 1'b0;
assign COL[12396] = 1'b0;
assign COL[12397] = 1'b0;
assign COL[12398] = 1'b0;
assign COL[12399] = 1'b0;
assign COL[12400] = 1'b0;
assign COL[12401] = 1'b0;
assign COL[12402] = 1'b0;
assign COL[12403] = 1'b0;
assign COL[12404] = 1'b0;
assign COL[12405] = 1'b0;
assign COL[12406] = 1'b0;
assign COL[12407] = 1'b0;
assign COL[12408] = 1'b0;
assign COL[12409] = 1'b0;
assign COL[12410] = 1'b1;
assign COL[12411] = 1'b1;
assign COL[12412] = 1'b1;
assign COL[12413] = 1'b1;
assign COL[12414] = 1'b1;
assign COL[12415] = 1'b0;
assign COL[12416] = 1'b0;
assign COL[12417] = 1'b0;
assign COL[12418] = 1'b0;
assign COL[12419] = 1'b0;
assign COL[12420] = 1'b0;
assign COL[12421] = 1'b0;
assign COL[12422] = 1'b0;
assign COL[12423] = 1'b0;
assign COL[12424] = 1'b0;
assign COL[12425] = 1'b0;
assign COL[12426] = 1'b0;
assign COL[12427] = 1'b0;
assign COL[12428] = 1'b0;
assign COL[12429] = 1'b0;
assign COL[12430] = 1'b0;
assign COL[12431] = 1'b0;
assign COL[12432] = 1'b0;
assign COL[12433] = 1'b0;
assign COL[12434] = 1'b0;
assign COL[12435] = 1'b0;
assign COL[12436] = 1'b0;
assign COL[12437] = 1'b0;
assign COL[12438] = 1'b0;
assign COL[12439] = 1'b0;
assign COL[12440] = 1'b0;
assign COL[12441] = 1'b0;
assign COL[12442] = 1'b0;
assign COL[12443] = 1'b0;
assign COL[12444] = 1'b0;
assign COL[12445] = 1'b0;
assign COL[12446] = 1'b0;
assign COL[12447] = 1'b0;
assign COL[12448] = 1'b0;
assign COL[12449] = 1'b0;
assign COL[12450] = 1'b0;
assign COL[12451] = 1'b0;
assign COL[12452] = 1'b0;
assign COL[12453] = 1'b0;
assign COL[12454] = 1'b0;
assign COL[12455] = 1'b0;
assign COL[12456] = 1'b0;
assign COL[12457] = 1'b0;
assign COL[12458] = 1'b0;
assign COL[12459] = 1'b0;
assign COL[12460] = 1'b0;
assign COL[12461] = 1'b0;
assign COL[12462] = 1'b0;
assign COL[12463] = 1'b0;
assign COL[12464] = 1'b0;
assign COL[12465] = 1'b0;
assign COL[12466] = 1'b0;
assign COL[12467] = 1'b0;
assign COL[12468] = 1'b0;
assign COL[12469] = 1'b0;
assign COL[12470] = 1'b0;
assign COL[12471] = 1'b0;
assign COL[12472] = 1'b0;
assign COL[12473] = 1'b0;
assign COL[12474] = 1'b0;
assign COL[12475] = 1'b0;
assign COL[12476] = 1'b0;
assign COL[12477] = 1'b0;
assign COL[12478] = 1'b0;
assign COL[12479] = 1'b0;
assign COL[12480] = 1'b0;
assign COL[12481] = 1'b1;
assign COL[12482] = 1'b1;
assign COL[12483] = 1'b1;
assign COL[12484] = 1'b1;
assign COL[12485] = 1'b0;
assign COL[12486] = 1'b0;
assign COL[12487] = 1'b0;
assign COL[12488] = 1'b0;
assign COL[12489] = 1'b0;
assign COL[12490] = 1'b0;
assign COL[12491] = 1'b1;
assign COL[12492] = 1'b1;
assign COL[12493] = 1'b1;
assign COL[12494] = 1'b1;
assign COL[12495] = 1'b1;
assign COL[12496] = 1'b1;
assign COL[12497] = 1'b1;
assign COL[12498] = 1'b1;
assign COL[12499] = 1'b1;
assign COL[12500] = 1'b1;
assign COL[12501] = 1'b1;
assign COL[12502] = 1'b1;
assign COL[12503] = 1'b1;
assign COL[12504] = 1'b1;
assign COL[12505] = 1'b1;
assign COL[12506] = 1'b1;
assign COL[12507] = 1'b1;
assign COL[12508] = 1'b1;
assign COL[12509] = 1'b1;
assign COL[12510] = 1'b1;
assign COL[12511] = 1'b1;
assign COL[12512] = 1'b1;
assign COL[12513] = 1'b1;
assign COL[12514] = 1'b1;
assign COL[12515] = 1'b1;
assign COL[12516] = 1'b1;
assign COL[12517] = 1'b1;
assign COL[12518] = 1'b1;
assign COL[12519] = 1'b1;
assign COL[12520] = 1'b1;
assign COL[12521] = 1'b1;
assign COL[12522] = 1'b1;
assign COL[12523] = 1'b1;
assign COL[12524] = 1'b1;
assign COL[12525] = 1'b1;
assign COL[12526] = 1'b1;
assign COL[12527] = 1'b1;
assign COL[12528] = 1'b1;
assign COL[12529] = 1'b0;
assign COL[12530] = 1'b0;
assign COL[12531] = 1'b0;
assign COL[12532] = 1'b0;
assign COL[12533] = 1'b0;
assign COL[12534] = 1'b0;
assign COL[12535] = 1'b1;
assign COL[12536] = 1'b1;
assign COL[12537] = 1'b1;
assign COL[12538] = 1'b1;
assign COL[12539] = 1'b0;
assign COL[12540] = 1'b0;
assign COL[12541] = 1'b0;
assign COL[12542] = 1'b0;
assign COL[12543] = 1'b0;
assign COL[12544] = 1'b0;
assign COL[12545] = 1'b0;
assign COL[12546] = 1'b0;
assign COL[12547] = 1'b0;
assign COL[12548] = 1'b0;
assign COL[12549] = 1'b0;
assign COL[12550] = 1'b0;
assign COL[12551] = 1'b0;
assign COL[12552] = 1'b0;
assign COL[12553] = 1'b0;
assign COL[12554] = 1'b0;
assign COL[12555] = 1'b0;
assign COL[12556] = 1'b0;
assign COL[12557] = 1'b0;
assign COL[12558] = 1'b0;
assign COL[12559] = 1'b0;
assign COL[12560] = 1'b0;
assign COL[12561] = 1'b0;
assign COL[12562] = 1'b0;
assign COL[12563] = 1'b0;
assign COL[12564] = 1'b0;
assign COL[12565] = 1'b0;
assign COL[12566] = 1'b0;
assign COL[12567] = 1'b0;
assign COL[12568] = 1'b0;
assign COL[12569] = 1'b0;
assign COL[12570] = 1'b1;
assign COL[12571] = 1'b1;
assign COL[12572] = 1'b1;
assign COL[12573] = 1'b1;
assign COL[12574] = 1'b1;
assign COL[12575] = 1'b0;
assign COL[12576] = 1'b0;
assign COL[12577] = 1'b0;
assign COL[12578] = 1'b0;
assign COL[12579] = 1'b0;
assign COL[12580] = 1'b0;
assign COL[12581] = 1'b0;
assign COL[12582] = 1'b0;
assign COL[12583] = 1'b0;
assign COL[12584] = 1'b0;
assign COL[12585] = 1'b0;
assign COL[12586] = 1'b0;
assign COL[12587] = 1'b0;
assign COL[12588] = 1'b0;
assign COL[12589] = 1'b0;
assign COL[12590] = 1'b0;
assign COL[12591] = 1'b0;
assign COL[12592] = 1'b0;
assign COL[12593] = 1'b0;
assign COL[12594] = 1'b0;
assign COL[12595] = 1'b0;
assign COL[12596] = 1'b0;
assign COL[12597] = 1'b0;
assign COL[12598] = 1'b0;
assign COL[12599] = 1'b0;
assign COL[12600] = 1'b0;
assign COL[12601] = 1'b0;
assign COL[12602] = 1'b0;
assign COL[12603] = 1'b0;
assign COL[12604] = 1'b0;
assign COL[12605] = 1'b0;
assign COL[12606] = 1'b0;
assign COL[12607] = 1'b0;
assign COL[12608] = 1'b0;
assign COL[12609] = 1'b0;
assign COL[12610] = 1'b0;
assign COL[12611] = 1'b0;
assign COL[12612] = 1'b0;
assign COL[12613] = 1'b0;
assign COL[12614] = 1'b0;
assign COL[12615] = 1'b0;
assign COL[12616] = 1'b0;
assign COL[12617] = 1'b0;
assign COL[12618] = 1'b0;
assign COL[12619] = 1'b0;
assign COL[12620] = 1'b0;
assign COL[12621] = 1'b0;
assign COL[12622] = 1'b0;
assign COL[12623] = 1'b0;
assign COL[12624] = 1'b0;
assign COL[12625] = 1'b0;
assign COL[12626] = 1'b0;
assign COL[12627] = 1'b0;
assign COL[12628] = 1'b0;
assign COL[12629] = 1'b0;
assign COL[12630] = 1'b0;
assign COL[12631] = 1'b0;
assign COL[12632] = 1'b0;
assign COL[12633] = 1'b0;
assign COL[12634] = 1'b0;
assign COL[12635] = 1'b0;
assign COL[12636] = 1'b0;
assign COL[12637] = 1'b0;
assign COL[12638] = 1'b0;
assign COL[12639] = 1'b0;
assign COL[12640] = 1'b0;
assign COL[12641] = 1'b1;
assign COL[12642] = 1'b1;
assign COL[12643] = 1'b1;
assign COL[12644] = 1'b1;
assign COL[12645] = 1'b0;
assign COL[12646] = 1'b0;
assign COL[12647] = 1'b0;
assign COL[12648] = 1'b0;
assign COL[12649] = 1'b0;
assign COL[12650] = 1'b0;
assign COL[12651] = 1'b1;
assign COL[12652] = 1'b1;
assign COL[12653] = 1'b1;
assign COL[12654] = 1'b1;
assign COL[12655] = 1'b1;
assign COL[12656] = 1'b1;
assign COL[12657] = 1'b1;
assign COL[12658] = 1'b1;
assign COL[12659] = 1'b1;
assign COL[12660] = 1'b1;
assign COL[12661] = 1'b1;
assign COL[12662] = 1'b1;
assign COL[12663] = 1'b1;
assign COL[12664] = 1'b1;
assign COL[12665] = 1'b1;
assign COL[12666] = 1'b1;
assign COL[12667] = 1'b1;
assign COL[12668] = 1'b1;
assign COL[12669] = 1'b1;
assign COL[12670] = 1'b1;
assign COL[12671] = 1'b1;
assign COL[12672] = 1'b1;
assign COL[12673] = 1'b1;
assign COL[12674] = 1'b1;
assign COL[12675] = 1'b1;
assign COL[12676] = 1'b1;
assign COL[12677] = 1'b1;
assign COL[12678] = 1'b1;
assign COL[12679] = 1'b1;
assign COL[12680] = 1'b1;
assign COL[12681] = 1'b1;
assign COL[12682] = 1'b1;
assign COL[12683] = 1'b1;
assign COL[12684] = 1'b1;
assign COL[12685] = 1'b1;
assign COL[12686] = 1'b1;
assign COL[12687] = 1'b1;
assign COL[12688] = 1'b1;
assign COL[12689] = 1'b0;
assign COL[12690] = 1'b0;
assign COL[12691] = 1'b0;
assign COL[12692] = 1'b0;
assign COL[12693] = 1'b0;
assign COL[12694] = 1'b0;
assign COL[12695] = 1'b1;
assign COL[12696] = 1'b1;
assign COL[12697] = 1'b1;
assign COL[12698] = 1'b1;
assign COL[12699] = 1'b0;
assign COL[12700] = 1'b0;
assign COL[12701] = 1'b0;
assign COL[12702] = 1'b0;
assign COL[12703] = 1'b0;
assign COL[12704] = 1'b0;
assign COL[12705] = 1'b0;
assign COL[12706] = 1'b0;
assign COL[12707] = 1'b0;
assign COL[12708] = 1'b0;
assign COL[12709] = 1'b0;
assign COL[12710] = 1'b0;
assign COL[12711] = 1'b0;
assign COL[12712] = 1'b0;
assign COL[12713] = 1'b0;
assign COL[12714] = 1'b0;
assign COL[12715] = 1'b0;
assign COL[12716] = 1'b0;
assign COL[12717] = 1'b0;
assign COL[12718] = 1'b0;
assign COL[12719] = 1'b0;
assign COL[12720] = 1'b0;
assign COL[12721] = 1'b0;
assign COL[12722] = 1'b0;
assign COL[12723] = 1'b0;
assign COL[12724] = 1'b0;
assign COL[12725] = 1'b0;
assign COL[12726] = 1'b0;
assign COL[12727] = 1'b0;
assign COL[12728] = 1'b0;
assign COL[12729] = 1'b0;
assign COL[12730] = 1'b1;
assign COL[12731] = 1'b1;
assign COL[12732] = 1'b1;
assign COL[12733] = 1'b1;
assign COL[12734] = 1'b1;
assign COL[12735] = 1'b0;
assign COL[12736] = 1'b0;
assign COL[12737] = 1'b0;
assign COL[12738] = 1'b0;
assign COL[12739] = 1'b0;
assign COL[12740] = 1'b0;
assign COL[12741] = 1'b0;
assign COL[12742] = 1'b0;
assign COL[12743] = 1'b0;
assign COL[12744] = 1'b0;
assign COL[12745] = 1'b0;
assign COL[12746] = 1'b0;
assign COL[12747] = 1'b0;
assign COL[12748] = 1'b0;
assign COL[12749] = 1'b0;
assign COL[12750] = 1'b0;
assign COL[12751] = 1'b0;
assign COL[12752] = 1'b0;
assign COL[12753] = 1'b0;
assign COL[12754] = 1'b0;
assign COL[12755] = 1'b0;
assign COL[12756] = 1'b0;
assign COL[12757] = 1'b0;
assign COL[12758] = 1'b0;
assign COL[12759] = 1'b0;
assign COL[12760] = 1'b0;
assign COL[12761] = 1'b0;
assign COL[12762] = 1'b0;
assign COL[12763] = 1'b0;
assign COL[12764] = 1'b0;
assign COL[12765] = 1'b0;
assign COL[12766] = 1'b0;
assign COL[12767] = 1'b0;
assign COL[12768] = 1'b0;
assign COL[12769] = 1'b0;
assign COL[12770] = 1'b0;
assign COL[12771] = 1'b0;
assign COL[12772] = 1'b0;
assign COL[12773] = 1'b0;
assign COL[12774] = 1'b0;
assign COL[12775] = 1'b0;
assign COL[12776] = 1'b0;
assign COL[12777] = 1'b0;
assign COL[12778] = 1'b0;
assign COL[12779] = 1'b0;
assign COL[12780] = 1'b0;
assign COL[12781] = 1'b0;
assign COL[12782] = 1'b0;
assign COL[12783] = 1'b0;
assign COL[12784] = 1'b0;
assign COL[12785] = 1'b0;
assign COL[12786] = 1'b0;
assign COL[12787] = 1'b0;
assign COL[12788] = 1'b0;
assign COL[12789] = 1'b0;
assign COL[12790] = 1'b0;
assign COL[12791] = 1'b0;
assign COL[12792] = 1'b0;
assign COL[12793] = 1'b0;
assign COL[12794] = 1'b0;
assign COL[12795] = 1'b0;
assign COL[12796] = 1'b0;
assign COL[12797] = 1'b0;
assign COL[12798] = 1'b0;
assign COL[12799] = 1'b0;
assign COL[12800] = 1'b0;
assign COL[12801] = 1'b1;
assign COL[12802] = 1'b1;
assign COL[12803] = 1'b1;
assign COL[12804] = 1'b1;
assign COL[12805] = 1'b0;
assign COL[12806] = 1'b0;
assign COL[12807] = 1'b0;
assign COL[12808] = 1'b0;
assign COL[12809] = 1'b0;
assign COL[12810] = 1'b0;
assign COL[12811] = 1'b1;
assign COL[12812] = 1'b1;
assign COL[12813] = 1'b1;
assign COL[12814] = 1'b1;
assign COL[12815] = 1'b1;
assign COL[12816] = 1'b1;
assign COL[12817] = 1'b1;
assign COL[12818] = 1'b1;
assign COL[12819] = 1'b1;
assign COL[12820] = 1'b1;
assign COL[12821] = 1'b1;
assign COL[12822] = 1'b1;
assign COL[12823] = 1'b1;
assign COL[12824] = 1'b1;
assign COL[12825] = 1'b1;
assign COL[12826] = 1'b1;
assign COL[12827] = 1'b1;
assign COL[12828] = 1'b1;
assign COL[12829] = 1'b1;
assign COL[12830] = 1'b1;
assign COL[12831] = 1'b1;
assign COL[12832] = 1'b1;
assign COL[12833] = 1'b1;
assign COL[12834] = 1'b1;
assign COL[12835] = 1'b1;
assign COL[12836] = 1'b1;
assign COL[12837] = 1'b1;
assign COL[12838] = 1'b1;
assign COL[12839] = 1'b1;
assign COL[12840] = 1'b1;
assign COL[12841] = 1'b1;
assign COL[12842] = 1'b1;
assign COL[12843] = 1'b1;
assign COL[12844] = 1'b1;
assign COL[12845] = 1'b1;
assign COL[12846] = 1'b1;
assign COL[12847] = 1'b1;
assign COL[12848] = 1'b1;
assign COL[12849] = 1'b0;
assign COL[12850] = 1'b0;
assign COL[12851] = 1'b0;
assign COL[12852] = 1'b0;
assign COL[12853] = 1'b0;
assign COL[12854] = 1'b0;
assign COL[12855] = 1'b1;
assign COL[12856] = 1'b1;
assign COL[12857] = 1'b1;
assign COL[12858] = 1'b1;
assign COL[12859] = 1'b0;
assign COL[12860] = 1'b0;
assign COL[12861] = 1'b0;
assign COL[12862] = 1'b0;
assign COL[12863] = 1'b0;
assign COL[12864] = 1'b0;
assign COL[12865] = 1'b0;
assign COL[12866] = 1'b0;
assign COL[12867] = 1'b0;
assign COL[12868] = 1'b0;
assign COL[12869] = 1'b0;
assign COL[12870] = 1'b0;
assign COL[12871] = 1'b0;
assign COL[12872] = 1'b0;
assign COL[12873] = 1'b0;
assign COL[12874] = 1'b0;
assign COL[12875] = 1'b0;
assign COL[12876] = 1'b0;
assign COL[12877] = 1'b0;
assign COL[12878] = 1'b0;
assign COL[12879] = 1'b0;
assign COL[12880] = 1'b0;
assign COL[12881] = 1'b0;
assign COL[12882] = 1'b0;
assign COL[12883] = 1'b0;
assign COL[12884] = 1'b0;
assign COL[12885] = 1'b0;
assign COL[12886] = 1'b0;
assign COL[12887] = 1'b0;
assign COL[12888] = 1'b0;
assign COL[12889] = 1'b0;
assign COL[12890] = 1'b1;
assign COL[12891] = 1'b1;
assign COL[12892] = 1'b1;
assign COL[12893] = 1'b1;
assign COL[12894] = 1'b1;
assign COL[12895] = 1'b0;
assign COL[12896] = 1'b0;
assign COL[12897] = 1'b0;
assign COL[12898] = 1'b0;
assign COL[12899] = 1'b0;
assign COL[12900] = 1'b0;
assign COL[12901] = 1'b0;
assign COL[12902] = 1'b0;
assign COL[12903] = 1'b0;
assign COL[12904] = 1'b0;
assign COL[12905] = 1'b0;
assign COL[12906] = 1'b0;
assign COL[12907] = 1'b0;
assign COL[12908] = 1'b0;
assign COL[12909] = 1'b0;
assign COL[12910] = 1'b0;
assign COL[12911] = 1'b0;
assign COL[12912] = 1'b0;
assign COL[12913] = 1'b0;
assign COL[12914] = 1'b0;
assign COL[12915] = 1'b0;
assign COL[12916] = 1'b0;
assign COL[12917] = 1'b0;
assign COL[12918] = 1'b0;
assign COL[12919] = 1'b0;
assign COL[12920] = 1'b0;
assign COL[12921] = 1'b0;
assign COL[12922] = 1'b0;
assign COL[12923] = 1'b0;
assign COL[12924] = 1'b0;
assign COL[12925] = 1'b0;
assign COL[12926] = 1'b0;
assign COL[12927] = 1'b0;
assign COL[12928] = 1'b0;
assign COL[12929] = 1'b0;
assign COL[12930] = 1'b0;
assign COL[12931] = 1'b0;
assign COL[12932] = 1'b0;
assign COL[12933] = 1'b0;
assign COL[12934] = 1'b0;
assign COL[12935] = 1'b0;
assign COL[12936] = 1'b0;
assign COL[12937] = 1'b0;
assign COL[12938] = 1'b0;
assign COL[12939] = 1'b0;
assign COL[12940] = 1'b0;
assign COL[12941] = 1'b0;
assign COL[12942] = 1'b0;
assign COL[12943] = 1'b0;
assign COL[12944] = 1'b0;
assign COL[12945] = 1'b0;
assign COL[12946] = 1'b0;
assign COL[12947] = 1'b0;
assign COL[12948] = 1'b0;
assign COL[12949] = 1'b0;
assign COL[12950] = 1'b0;
assign COL[12951] = 1'b0;
assign COL[12952] = 1'b0;
assign COL[12953] = 1'b0;
assign COL[12954] = 1'b0;
assign COL[12955] = 1'b0;
assign COL[12956] = 1'b0;
assign COL[12957] = 1'b0;
assign COL[12958] = 1'b0;
assign COL[12959] = 1'b0;
assign COL[12960] = 1'b0;
assign COL[12961] = 1'b1;
assign COL[12962] = 1'b1;
assign COL[12963] = 1'b1;
assign COL[12964] = 1'b1;
assign COL[12965] = 1'b0;
assign COL[12966] = 1'b0;
assign COL[12967] = 1'b0;
assign COL[12968] = 1'b0;
assign COL[12969] = 1'b0;
assign COL[12970] = 1'b0;
assign COL[12971] = 1'b0;
assign COL[12972] = 1'b0;
assign COL[12973] = 1'b0;
assign COL[12974] = 1'b0;
assign COL[12975] = 1'b0;
assign COL[12976] = 1'b0;
assign COL[12977] = 1'b0;
assign COL[12978] = 1'b0;
assign COL[12979] = 1'b0;
assign COL[12980] = 1'b0;
assign COL[12981] = 1'b0;
assign COL[12982] = 1'b0;
assign COL[12983] = 1'b0;
assign COL[12984] = 1'b0;
assign COL[12985] = 1'b0;
assign COL[12986] = 1'b0;
assign COL[12987] = 1'b0;
assign COL[12988] = 1'b0;
assign COL[12989] = 1'b0;
assign COL[12990] = 1'b0;
assign COL[12991] = 1'b0;
assign COL[12992] = 1'b0;
assign COL[12993] = 1'b0;
assign COL[12994] = 1'b0;
assign COL[12995] = 1'b0;
assign COL[12996] = 1'b0;
assign COL[12997] = 1'b0;
assign COL[12998] = 1'b0;
assign COL[12999] = 1'b0;
assign COL[13000] = 1'b0;
assign COL[13001] = 1'b0;
assign COL[13002] = 1'b0;
assign COL[13003] = 1'b0;
assign COL[13004] = 1'b0;
assign COL[13005] = 1'b0;
assign COL[13006] = 1'b0;
assign COL[13007] = 1'b0;
assign COL[13008] = 1'b0;
assign COL[13009] = 1'b0;
assign COL[13010] = 1'b0;
assign COL[13011] = 1'b0;
assign COL[13012] = 1'b0;
assign COL[13013] = 1'b0;
assign COL[13014] = 1'b0;
assign COL[13015] = 1'b1;
assign COL[13016] = 1'b1;
assign COL[13017] = 1'b1;
assign COL[13018] = 1'b1;
assign COL[13019] = 1'b0;
assign COL[13020] = 1'b0;
assign COL[13021] = 1'b0;
assign COL[13022] = 1'b0;
assign COL[13023] = 1'b0;
assign COL[13024] = 1'b0;
assign COL[13025] = 1'b0;
assign COL[13026] = 1'b0;
assign COL[13027] = 1'b0;
assign COL[13028] = 1'b0;
assign COL[13029] = 1'b0;
assign COL[13030] = 1'b0;
assign COL[13031] = 1'b0;
assign COL[13032] = 1'b0;
assign COL[13033] = 1'b0;
assign COL[13034] = 1'b0;
assign COL[13035] = 1'b0;
assign COL[13036] = 1'b0;
assign COL[13037] = 1'b0;
assign COL[13038] = 1'b0;
assign COL[13039] = 1'b0;
assign COL[13040] = 1'b0;
assign COL[13041] = 1'b0;
assign COL[13042] = 1'b0;
assign COL[13043] = 1'b0;
assign COL[13044] = 1'b0;
assign COL[13045] = 1'b0;
assign COL[13046] = 1'b0;
assign COL[13047] = 1'b0;
assign COL[13048] = 1'b0;
assign COL[13049] = 1'b0;
assign COL[13050] = 1'b1;
assign COL[13051] = 1'b1;
assign COL[13052] = 1'b1;
assign COL[13053] = 1'b1;
assign COL[13054] = 1'b1;
assign COL[13055] = 1'b0;
assign COL[13056] = 1'b0;
assign COL[13057] = 1'b0;
assign COL[13058] = 1'b0;
assign COL[13059] = 1'b0;
assign COL[13060] = 1'b0;
assign COL[13061] = 1'b0;
assign COL[13062] = 1'b0;
assign COL[13063] = 1'b0;
assign COL[13064] = 1'b0;
assign COL[13065] = 1'b0;
assign COL[13066] = 1'b0;
assign COL[13067] = 1'b0;
assign COL[13068] = 1'b0;
assign COL[13069] = 1'b0;
assign COL[13070] = 1'b0;
assign COL[13071] = 1'b0;
assign COL[13072] = 1'b0;
assign COL[13073] = 1'b0;
assign COL[13074] = 1'b0;
assign COL[13075] = 1'b0;
assign COL[13076] = 1'b0;
assign COL[13077] = 1'b0;
assign COL[13078] = 1'b0;
assign COL[13079] = 1'b0;
assign COL[13080] = 1'b0;
assign COL[13081] = 1'b0;
assign COL[13082] = 1'b0;
assign COL[13083] = 1'b0;
assign COL[13084] = 1'b0;
assign COL[13085] = 1'b0;
assign COL[13086] = 1'b0;
assign COL[13087] = 1'b0;
assign COL[13088] = 1'b0;
assign COL[13089] = 1'b0;
assign COL[13090] = 1'b0;
assign COL[13091] = 1'b0;
assign COL[13092] = 1'b0;
assign COL[13093] = 1'b0;
assign COL[13094] = 1'b0;
assign COL[13095] = 1'b0;
assign COL[13096] = 1'b0;
assign COL[13097] = 1'b0;
assign COL[13098] = 1'b0;
assign COL[13099] = 1'b0;
assign COL[13100] = 1'b0;
assign COL[13101] = 1'b0;
assign COL[13102] = 1'b0;
assign COL[13103] = 1'b0;
assign COL[13104] = 1'b0;
assign COL[13105] = 1'b0;
assign COL[13106] = 1'b0;
assign COL[13107] = 1'b0;
assign COL[13108] = 1'b0;
assign COL[13109] = 1'b0;
assign COL[13110] = 1'b0;
assign COL[13111] = 1'b0;
assign COL[13112] = 1'b0;
assign COL[13113] = 1'b0;
assign COL[13114] = 1'b0;
assign COL[13115] = 1'b0;
assign COL[13116] = 1'b0;
assign COL[13117] = 1'b0;
assign COL[13118] = 1'b0;
assign COL[13119] = 1'b0;
assign COL[13120] = 1'b0;
assign COL[13121] = 1'b1;
assign COL[13122] = 1'b1;
assign COL[13123] = 1'b1;
assign COL[13124] = 1'b1;
assign COL[13125] = 1'b0;
assign COL[13126] = 1'b0;
assign COL[13127] = 1'b0;
assign COL[13128] = 1'b0;
assign COL[13129] = 1'b0;
assign COL[13130] = 1'b0;
assign COL[13131] = 1'b0;
assign COL[13132] = 1'b0;
assign COL[13133] = 1'b0;
assign COL[13134] = 1'b0;
assign COL[13135] = 1'b0;
assign COL[13136] = 1'b0;
assign COL[13137] = 1'b0;
assign COL[13138] = 1'b0;
assign COL[13139] = 1'b0;
assign COL[13140] = 1'b0;
assign COL[13141] = 1'b0;
assign COL[13142] = 1'b0;
assign COL[13143] = 1'b0;
assign COL[13144] = 1'b0;
assign COL[13145] = 1'b0;
assign COL[13146] = 1'b0;
assign COL[13147] = 1'b0;
assign COL[13148] = 1'b0;
assign COL[13149] = 1'b0;
assign COL[13150] = 1'b0;
assign COL[13151] = 1'b0;
assign COL[13152] = 1'b0;
assign COL[13153] = 1'b0;
assign COL[13154] = 1'b0;
assign COL[13155] = 1'b0;
assign COL[13156] = 1'b0;
assign COL[13157] = 1'b0;
assign COL[13158] = 1'b0;
assign COL[13159] = 1'b0;
assign COL[13160] = 1'b0;
assign COL[13161] = 1'b0;
assign COL[13162] = 1'b0;
assign COL[13163] = 1'b0;
assign COL[13164] = 1'b0;
assign COL[13165] = 1'b0;
assign COL[13166] = 1'b0;
assign COL[13167] = 1'b0;
assign COL[13168] = 1'b0;
assign COL[13169] = 1'b0;
assign COL[13170] = 1'b0;
assign COL[13171] = 1'b0;
assign COL[13172] = 1'b0;
assign COL[13173] = 1'b0;
assign COL[13174] = 1'b0;
assign COL[13175] = 1'b1;
assign COL[13176] = 1'b1;
assign COL[13177] = 1'b1;
assign COL[13178] = 1'b1;
assign COL[13179] = 1'b0;
assign COL[13180] = 1'b0;
assign COL[13181] = 1'b0;
assign COL[13182] = 1'b0;
assign COL[13183] = 1'b0;
assign COL[13184] = 1'b0;
assign COL[13185] = 1'b0;
assign COL[13186] = 1'b0;
assign COL[13187] = 1'b0;
assign COL[13188] = 1'b0;
assign COL[13189] = 1'b0;
assign COL[13190] = 1'b0;
assign COL[13191] = 1'b0;
assign COL[13192] = 1'b0;
assign COL[13193] = 1'b0;
assign COL[13194] = 1'b0;
assign COL[13195] = 1'b0;
assign COL[13196] = 1'b0;
assign COL[13197] = 1'b0;
assign COL[13198] = 1'b0;
assign COL[13199] = 1'b0;
assign COL[13200] = 1'b0;
assign COL[13201] = 1'b0;
assign COL[13202] = 1'b0;
assign COL[13203] = 1'b0;
assign COL[13204] = 1'b0;
assign COL[13205] = 1'b0;
assign COL[13206] = 1'b0;
assign COL[13207] = 1'b0;
assign COL[13208] = 1'b0;
assign COL[13209] = 1'b0;
assign COL[13210] = 1'b1;
assign COL[13211] = 1'b1;
assign COL[13212] = 1'b1;
assign COL[13213] = 1'b1;
assign COL[13214] = 1'b1;
assign COL[13215] = 1'b0;
assign COL[13216] = 1'b0;
assign COL[13217] = 1'b0;
assign COL[13218] = 1'b0;
assign COL[13219] = 1'b0;
assign COL[13220] = 1'b0;
assign COL[13221] = 1'b0;
assign COL[13222] = 1'b0;
assign COL[13223] = 1'b0;
assign COL[13224] = 1'b0;
assign COL[13225] = 1'b0;
assign COL[13226] = 1'b0;
assign COL[13227] = 1'b0;
assign COL[13228] = 1'b0;
assign COL[13229] = 1'b0;
assign COL[13230] = 1'b0;
assign COL[13231] = 1'b0;
assign COL[13232] = 1'b0;
assign COL[13233] = 1'b0;
assign COL[13234] = 1'b0;
assign COL[13235] = 1'b0;
assign COL[13236] = 1'b0;
assign COL[13237] = 1'b0;
assign COL[13238] = 1'b0;
assign COL[13239] = 1'b0;
assign COL[13240] = 1'b0;
assign COL[13241] = 1'b0;
assign COL[13242] = 1'b0;
assign COL[13243] = 1'b0;
assign COL[13244] = 1'b0;
assign COL[13245] = 1'b0;
assign COL[13246] = 1'b0;
assign COL[13247] = 1'b0;
assign COL[13248] = 1'b0;
assign COL[13249] = 1'b0;
assign COL[13250] = 1'b0;
assign COL[13251] = 1'b0;
assign COL[13252] = 1'b0;
assign COL[13253] = 1'b0;
assign COL[13254] = 1'b0;
assign COL[13255] = 1'b0;
assign COL[13256] = 1'b0;
assign COL[13257] = 1'b0;
assign COL[13258] = 1'b0;
assign COL[13259] = 1'b0;
assign COL[13260] = 1'b0;
assign COL[13261] = 1'b0;
assign COL[13262] = 1'b0;
assign COL[13263] = 1'b0;
assign COL[13264] = 1'b0;
assign COL[13265] = 1'b0;
assign COL[13266] = 1'b0;
assign COL[13267] = 1'b0;
assign COL[13268] = 1'b0;
assign COL[13269] = 1'b0;
assign COL[13270] = 1'b0;
assign COL[13271] = 1'b0;
assign COL[13272] = 1'b0;
assign COL[13273] = 1'b0;
assign COL[13274] = 1'b0;
assign COL[13275] = 1'b0;
assign COL[13276] = 1'b0;
assign COL[13277] = 1'b0;
assign COL[13278] = 1'b0;
assign COL[13279] = 1'b0;
assign COL[13280] = 1'b0;
assign COL[13281] = 1'b1;
assign COL[13282] = 1'b1;
assign COL[13283] = 1'b1;
assign COL[13284] = 1'b1;
assign COL[13285] = 1'b0;
assign COL[13286] = 1'b0;
assign COL[13287] = 1'b0;
assign COL[13288] = 1'b0;
assign COL[13289] = 1'b0;
assign COL[13290] = 1'b0;
assign COL[13291] = 1'b0;
assign COL[13292] = 1'b0;
assign COL[13293] = 1'b0;
assign COL[13294] = 1'b0;
assign COL[13295] = 1'b0;
assign COL[13296] = 1'b0;
assign COL[13297] = 1'b0;
assign COL[13298] = 1'b0;
assign COL[13299] = 1'b0;
assign COL[13300] = 1'b0;
assign COL[13301] = 1'b0;
assign COL[13302] = 1'b0;
assign COL[13303] = 1'b0;
assign COL[13304] = 1'b0;
assign COL[13305] = 1'b0;
assign COL[13306] = 1'b0;
assign COL[13307] = 1'b0;
assign COL[13308] = 1'b0;
assign COL[13309] = 1'b0;
assign COL[13310] = 1'b0;
assign COL[13311] = 1'b0;
assign COL[13312] = 1'b0;
assign COL[13313] = 1'b0;
assign COL[13314] = 1'b0;
assign COL[13315] = 1'b0;
assign COL[13316] = 1'b0;
assign COL[13317] = 1'b0;
assign COL[13318] = 1'b0;
assign COL[13319] = 1'b0;
assign COL[13320] = 1'b0;
assign COL[13321] = 1'b0;
assign COL[13322] = 1'b0;
assign COL[13323] = 1'b0;
assign COL[13324] = 1'b0;
assign COL[13325] = 1'b0;
assign COL[13326] = 1'b0;
assign COL[13327] = 1'b0;
assign COL[13328] = 1'b0;
assign COL[13329] = 1'b0;
assign COL[13330] = 1'b0;
assign COL[13331] = 1'b0;
assign COL[13332] = 1'b0;
assign COL[13333] = 1'b0;
assign COL[13334] = 1'b0;
assign COL[13335] = 1'b1;
assign COL[13336] = 1'b1;
assign COL[13337] = 1'b1;
assign COL[13338] = 1'b1;
assign COL[13339] = 1'b0;
assign COL[13340] = 1'b0;
assign COL[13341] = 1'b0;
assign COL[13342] = 1'b0;
assign COL[13343] = 1'b0;
assign COL[13344] = 1'b0;
assign COL[13345] = 1'b0;
assign COL[13346] = 1'b0;
assign COL[13347] = 1'b0;
assign COL[13348] = 1'b0;
assign COL[13349] = 1'b0;
assign COL[13350] = 1'b0;
assign COL[13351] = 1'b0;
assign COL[13352] = 1'b0;
assign COL[13353] = 1'b0;
assign COL[13354] = 1'b0;
assign COL[13355] = 1'b0;
assign COL[13356] = 1'b0;
assign COL[13357] = 1'b0;
assign COL[13358] = 1'b0;
assign COL[13359] = 1'b0;
assign COL[13360] = 1'b0;
assign COL[13361] = 1'b0;
assign COL[13362] = 1'b0;
assign COL[13363] = 1'b0;
assign COL[13364] = 1'b0;
assign COL[13365] = 1'b0;
assign COL[13366] = 1'b0;
assign COL[13367] = 1'b0;
assign COL[13368] = 1'b0;
assign COL[13369] = 1'b0;
assign COL[13370] = 1'b1;
assign COL[13371] = 1'b1;
assign COL[13372] = 1'b1;
assign COL[13373] = 1'b1;
assign COL[13374] = 1'b1;
assign COL[13375] = 1'b0;
assign COL[13376] = 1'b0;
assign COL[13377] = 1'b0;
assign COL[13378] = 1'b0;
assign COL[13379] = 1'b0;
assign COL[13380] = 1'b0;
assign COL[13381] = 1'b0;
assign COL[13382] = 1'b0;
assign COL[13383] = 1'b0;
assign COL[13384] = 1'b0;
assign COL[13385] = 1'b0;
assign COL[13386] = 1'b0;
assign COL[13387] = 1'b0;
assign COL[13388] = 1'b0;
assign COL[13389] = 1'b0;
assign COL[13390] = 1'b0;
assign COL[13391] = 1'b0;
assign COL[13392] = 1'b0;
assign COL[13393] = 1'b0;
assign COL[13394] = 1'b0;
assign COL[13395] = 1'b0;
assign COL[13396] = 1'b0;
assign COL[13397] = 1'b0;
assign COL[13398] = 1'b0;
assign COL[13399] = 1'b0;
assign COL[13400] = 1'b0;
assign COL[13401] = 1'b0;
assign COL[13402] = 1'b0;
assign COL[13403] = 1'b0;
assign COL[13404] = 1'b0;
assign COL[13405] = 1'b0;
assign COL[13406] = 1'b0;
assign COL[13407] = 1'b0;
assign COL[13408] = 1'b0;
assign COL[13409] = 1'b0;
assign COL[13410] = 1'b0;
assign COL[13411] = 1'b0;
assign COL[13412] = 1'b0;
assign COL[13413] = 1'b0;
assign COL[13414] = 1'b0;
assign COL[13415] = 1'b0;
assign COL[13416] = 1'b0;
assign COL[13417] = 1'b0;
assign COL[13418] = 1'b0;
assign COL[13419] = 1'b0;
assign COL[13420] = 1'b0;
assign COL[13421] = 1'b0;
assign COL[13422] = 1'b0;
assign COL[13423] = 1'b0;
assign COL[13424] = 1'b0;
assign COL[13425] = 1'b0;
assign COL[13426] = 1'b0;
assign COL[13427] = 1'b0;
assign COL[13428] = 1'b0;
assign COL[13429] = 1'b0;
assign COL[13430] = 1'b0;
assign COL[13431] = 1'b0;
assign COL[13432] = 1'b0;
assign COL[13433] = 1'b0;
assign COL[13434] = 1'b0;
assign COL[13435] = 1'b0;
assign COL[13436] = 1'b0;
assign COL[13437] = 1'b0;
assign COL[13438] = 1'b0;
assign COL[13439] = 1'b0;
assign COL[13440] = 1'b0;
assign COL[13441] = 1'b1;
assign COL[13442] = 1'b1;
assign COL[13443] = 1'b1;
assign COL[13444] = 1'b1;
assign COL[13445] = 1'b0;
assign COL[13446] = 1'b0;
assign COL[13447] = 1'b0;
assign COL[13448] = 1'b0;
assign COL[13449] = 1'b0;
assign COL[13450] = 1'b0;
assign COL[13451] = 1'b0;
assign COL[13452] = 1'b0;
assign COL[13453] = 1'b0;
assign COL[13454] = 1'b0;
assign COL[13455] = 1'b0;
assign COL[13456] = 1'b0;
assign COL[13457] = 1'b0;
assign COL[13458] = 1'b0;
assign COL[13459] = 1'b0;
assign COL[13460] = 1'b0;
assign COL[13461] = 1'b0;
assign COL[13462] = 1'b0;
assign COL[13463] = 1'b0;
assign COL[13464] = 1'b0;
assign COL[13465] = 1'b0;
assign COL[13466] = 1'b0;
assign COL[13467] = 1'b0;
assign COL[13468] = 1'b0;
assign COL[13469] = 1'b0;
assign COL[13470] = 1'b0;
assign COL[13471] = 1'b0;
assign COL[13472] = 1'b0;
assign COL[13473] = 1'b0;
assign COL[13474] = 1'b0;
assign COL[13475] = 1'b0;
assign COL[13476] = 1'b0;
assign COL[13477] = 1'b0;
assign COL[13478] = 1'b0;
assign COL[13479] = 1'b0;
assign COL[13480] = 1'b0;
assign COL[13481] = 1'b0;
assign COL[13482] = 1'b0;
assign COL[13483] = 1'b0;
assign COL[13484] = 1'b0;
assign COL[13485] = 1'b0;
assign COL[13486] = 1'b0;
assign COL[13487] = 1'b0;
assign COL[13488] = 1'b0;
assign COL[13489] = 1'b0;
assign COL[13490] = 1'b0;
assign COL[13491] = 1'b0;
assign COL[13492] = 1'b0;
assign COL[13493] = 1'b0;
assign COL[13494] = 1'b0;
assign COL[13495] = 1'b1;
assign COL[13496] = 1'b1;
assign COL[13497] = 1'b1;
assign COL[13498] = 1'b1;
assign COL[13499] = 1'b0;
assign COL[13500] = 1'b0;
assign COL[13501] = 1'b0;
assign COL[13502] = 1'b0;
assign COL[13503] = 1'b0;
assign COL[13504] = 1'b0;
assign COL[13505] = 1'b0;
assign COL[13506] = 1'b0;
assign COL[13507] = 1'b0;
assign COL[13508] = 1'b0;
assign COL[13509] = 1'b0;
assign COL[13510] = 1'b0;
assign COL[13511] = 1'b0;
assign COL[13512] = 1'b0;
assign COL[13513] = 1'b0;
assign COL[13514] = 1'b0;
assign COL[13515] = 1'b0;
assign COL[13516] = 1'b0;
assign COL[13517] = 1'b0;
assign COL[13518] = 1'b0;
assign COL[13519] = 1'b0;
assign COL[13520] = 1'b0;
assign COL[13521] = 1'b0;
assign COL[13522] = 1'b0;
assign COL[13523] = 1'b0;
assign COL[13524] = 1'b0;
assign COL[13525] = 1'b0;
assign COL[13526] = 1'b0;
assign COL[13527] = 1'b0;
assign COL[13528] = 1'b0;
assign COL[13529] = 1'b0;
assign COL[13530] = 1'b1;
assign COL[13531] = 1'b1;
assign COL[13532] = 1'b1;
assign COL[13533] = 1'b1;
assign COL[13534] = 1'b1;
assign COL[13535] = 1'b0;
assign COL[13536] = 1'b0;
assign COL[13537] = 1'b0;
assign COL[13538] = 1'b0;
assign COL[13539] = 1'b0;
assign COL[13540] = 1'b0;
assign COL[13541] = 1'b0;
assign COL[13542] = 1'b0;
assign COL[13543] = 1'b0;
assign COL[13544] = 1'b0;
assign COL[13545] = 1'b0;
assign COL[13546] = 1'b0;
assign COL[13547] = 1'b0;
assign COL[13548] = 1'b0;
assign COL[13549] = 1'b0;
assign COL[13550] = 1'b0;
assign COL[13551] = 1'b0;
assign COL[13552] = 1'b0;
assign COL[13553] = 1'b0;
assign COL[13554] = 1'b0;
assign COL[13555] = 1'b0;
assign COL[13556] = 1'b0;
assign COL[13557] = 1'b0;
assign COL[13558] = 1'b0;
assign COL[13559] = 1'b0;
assign COL[13560] = 1'b0;
assign COL[13561] = 1'b0;
assign COL[13562] = 1'b0;
assign COL[13563] = 1'b0;
assign COL[13564] = 1'b0;
assign COL[13565] = 1'b0;
assign COL[13566] = 1'b0;
assign COL[13567] = 1'b0;
assign COL[13568] = 1'b0;
assign COL[13569] = 1'b0;
assign COL[13570] = 1'b0;
assign COL[13571] = 1'b0;
assign COL[13572] = 1'b0;
assign COL[13573] = 1'b0;
assign COL[13574] = 1'b0;
assign COL[13575] = 1'b0;
assign COL[13576] = 1'b0;
assign COL[13577] = 1'b0;
assign COL[13578] = 1'b0;
assign COL[13579] = 1'b0;
assign COL[13580] = 1'b0;
assign COL[13581] = 1'b0;
assign COL[13582] = 1'b0;
assign COL[13583] = 1'b0;
assign COL[13584] = 1'b0;
assign COL[13585] = 1'b0;
assign COL[13586] = 1'b0;
assign COL[13587] = 1'b0;
assign COL[13588] = 1'b0;
assign COL[13589] = 1'b0;
assign COL[13590] = 1'b0;
assign COL[13591] = 1'b0;
assign COL[13592] = 1'b0;
assign COL[13593] = 1'b0;
assign COL[13594] = 1'b0;
assign COL[13595] = 1'b0;
assign COL[13596] = 1'b0;
assign COL[13597] = 1'b0;
assign COL[13598] = 1'b0;
assign COL[13599] = 1'b0;
assign COL[13600] = 1'b0;
assign COL[13601] = 1'b1;
assign COL[13602] = 1'b1;
assign COL[13603] = 1'b1;
assign COL[13604] = 1'b1;
assign COL[13605] = 1'b0;
assign COL[13606] = 1'b0;
assign COL[13607] = 1'b0;
assign COL[13608] = 1'b0;
assign COL[13609] = 1'b0;
assign COL[13610] = 1'b0;
assign COL[13611] = 1'b0;
assign COL[13612] = 1'b0;
assign COL[13613] = 1'b0;
assign COL[13614] = 1'b0;
assign COL[13615] = 1'b0;
assign COL[13616] = 1'b0;
assign COL[13617] = 1'b0;
assign COL[13618] = 1'b0;
assign COL[13619] = 1'b0;
assign COL[13620] = 1'b0;
assign COL[13621] = 1'b0;
assign COL[13622] = 1'b0;
assign COL[13623] = 1'b0;
assign COL[13624] = 1'b0;
assign COL[13625] = 1'b0;
assign COL[13626] = 1'b0;
assign COL[13627] = 1'b0;
assign COL[13628] = 1'b0;
assign COL[13629] = 1'b0;
assign COL[13630] = 1'b0;
assign COL[13631] = 1'b0;
assign COL[13632] = 1'b0;
assign COL[13633] = 1'b0;
assign COL[13634] = 1'b0;
assign COL[13635] = 1'b0;
assign COL[13636] = 1'b0;
assign COL[13637] = 1'b0;
assign COL[13638] = 1'b0;
assign COL[13639] = 1'b0;
assign COL[13640] = 1'b0;
assign COL[13641] = 1'b0;
assign COL[13642] = 1'b0;
assign COL[13643] = 1'b0;
assign COL[13644] = 1'b0;
assign COL[13645] = 1'b0;
assign COL[13646] = 1'b0;
assign COL[13647] = 1'b0;
assign COL[13648] = 1'b0;
assign COL[13649] = 1'b0;
assign COL[13650] = 1'b0;
assign COL[13651] = 1'b0;
assign COL[13652] = 1'b0;
assign COL[13653] = 1'b0;
assign COL[13654] = 1'b0;
assign COL[13655] = 1'b1;
assign COL[13656] = 1'b1;
assign COL[13657] = 1'b1;
assign COL[13658] = 1'b1;
assign COL[13659] = 1'b0;
assign COL[13660] = 1'b0;
assign COL[13661] = 1'b0;
assign COL[13662] = 1'b0;
assign COL[13663] = 1'b0;
assign COL[13664] = 1'b0;
assign COL[13665] = 1'b0;
assign COL[13666] = 1'b0;
assign COL[13667] = 1'b0;
assign COL[13668] = 1'b0;
assign COL[13669] = 1'b0;
assign COL[13670] = 1'b0;
assign COL[13671] = 1'b0;
assign COL[13672] = 1'b0;
assign COL[13673] = 1'b0;
assign COL[13674] = 1'b0;
assign COL[13675] = 1'b0;
assign COL[13676] = 1'b0;
assign COL[13677] = 1'b0;
assign COL[13678] = 1'b0;
assign COL[13679] = 1'b0;
assign COL[13680] = 1'b0;
assign COL[13681] = 1'b0;
assign COL[13682] = 1'b0;
assign COL[13683] = 1'b0;
assign COL[13684] = 1'b0;
assign COL[13685] = 1'b0;
assign COL[13686] = 1'b0;
assign COL[13687] = 1'b0;
assign COL[13688] = 1'b0;
assign COL[13689] = 1'b0;
assign COL[13690] = 1'b1;
assign COL[13691] = 1'b1;
assign COL[13692] = 1'b1;
assign COL[13693] = 1'b1;
assign COL[13694] = 1'b1;
assign COL[13695] = 1'b0;
assign COL[13696] = 1'b0;
assign COL[13697] = 1'b0;
assign COL[13698] = 1'b0;
assign COL[13699] = 1'b0;
assign COL[13700] = 1'b0;
assign COL[13701] = 1'b0;
assign COL[13702] = 1'b0;
assign COL[13703] = 1'b0;
assign COL[13704] = 1'b0;
assign COL[13705] = 1'b0;
assign COL[13706] = 1'b0;
assign COL[13707] = 1'b0;
assign COL[13708] = 1'b0;
assign COL[13709] = 1'b0;
assign COL[13710] = 1'b0;
assign COL[13711] = 1'b0;
assign COL[13712] = 1'b0;
assign COL[13713] = 1'b0;
assign COL[13714] = 1'b0;
assign COL[13715] = 1'b0;
assign COL[13716] = 1'b0;
assign COL[13717] = 1'b0;
assign COL[13718] = 1'b0;
assign COL[13719] = 1'b0;
assign COL[13720] = 1'b0;
assign COL[13721] = 1'b0;
assign COL[13722] = 1'b0;
assign COL[13723] = 1'b0;
assign COL[13724] = 1'b0;
assign COL[13725] = 1'b0;
assign COL[13726] = 1'b0;
assign COL[13727] = 1'b0;
assign COL[13728] = 1'b0;
assign COL[13729] = 1'b0;
assign COL[13730] = 1'b0;
assign COL[13731] = 1'b0;
assign COL[13732] = 1'b0;
assign COL[13733] = 1'b0;
assign COL[13734] = 1'b0;
assign COL[13735] = 1'b0;
assign COL[13736] = 1'b0;
assign COL[13737] = 1'b0;
assign COL[13738] = 1'b0;
assign COL[13739] = 1'b0;
assign COL[13740] = 1'b0;
assign COL[13741] = 1'b0;
assign COL[13742] = 1'b0;
assign COL[13743] = 1'b0;
assign COL[13744] = 1'b0;
assign COL[13745] = 1'b0;
assign COL[13746] = 1'b0;
assign COL[13747] = 1'b0;
assign COL[13748] = 1'b0;
assign COL[13749] = 1'b0;
assign COL[13750] = 1'b0;
assign COL[13751] = 1'b0;
assign COL[13752] = 1'b0;
assign COL[13753] = 1'b0;
assign COL[13754] = 1'b0;
assign COL[13755] = 1'b0;
assign COL[13756] = 1'b0;
assign COL[13757] = 1'b0;
assign COL[13758] = 1'b0;
assign COL[13759] = 1'b0;
assign COL[13760] = 1'b0;
assign COL[13761] = 1'b1;
assign COL[13762] = 1'b1;
assign COL[13763] = 1'b1;
assign COL[13764] = 1'b1;
assign COL[13765] = 1'b0;
assign COL[13766] = 1'b0;
assign COL[13767] = 1'b0;
assign COL[13768] = 1'b0;
assign COL[13769] = 1'b0;
assign COL[13770] = 1'b0;
assign COL[13771] = 1'b0;
assign COL[13772] = 1'b0;
assign COL[13773] = 1'b0;
assign COL[13774] = 1'b0;
assign COL[13775] = 1'b0;
assign COL[13776] = 1'b0;
assign COL[13777] = 1'b0;
assign COL[13778] = 1'b0;
assign COL[13779] = 1'b0;
assign COL[13780] = 1'b0;
assign COL[13781] = 1'b0;
assign COL[13782] = 1'b0;
assign COL[13783] = 1'b0;
assign COL[13784] = 1'b0;
assign COL[13785] = 1'b0;
assign COL[13786] = 1'b0;
assign COL[13787] = 1'b0;
assign COL[13788] = 1'b0;
assign COL[13789] = 1'b0;
assign COL[13790] = 1'b0;
assign COL[13791] = 1'b0;
assign COL[13792] = 1'b0;
assign COL[13793] = 1'b0;
assign COL[13794] = 1'b0;
assign COL[13795] = 1'b0;
assign COL[13796] = 1'b0;
assign COL[13797] = 1'b0;
assign COL[13798] = 1'b0;
assign COL[13799] = 1'b0;
assign COL[13800] = 1'b0;
assign COL[13801] = 1'b0;
assign COL[13802] = 1'b0;
assign COL[13803] = 1'b0;
assign COL[13804] = 1'b0;
assign COL[13805] = 1'b0;
assign COL[13806] = 1'b0;
assign COL[13807] = 1'b0;
assign COL[13808] = 1'b0;
assign COL[13809] = 1'b0;
assign COL[13810] = 1'b0;
assign COL[13811] = 1'b0;
assign COL[13812] = 1'b0;
assign COL[13813] = 1'b0;
assign COL[13814] = 1'b0;
assign COL[13815] = 1'b1;
assign COL[13816] = 1'b1;
assign COL[13817] = 1'b1;
assign COL[13818] = 1'b1;
assign COL[13819] = 1'b0;
assign COL[13820] = 1'b0;
assign COL[13821] = 1'b0;
assign COL[13822] = 1'b0;
assign COL[13823] = 1'b0;
assign COL[13824] = 1'b0;
assign COL[13825] = 1'b0;
assign COL[13826] = 1'b0;
assign COL[13827] = 1'b0;
assign COL[13828] = 1'b0;
assign COL[13829] = 1'b0;
assign COL[13830] = 1'b0;
assign COL[13831] = 1'b0;
assign COL[13832] = 1'b0;
assign COL[13833] = 1'b0;
assign COL[13834] = 1'b0;
assign COL[13835] = 1'b0;
assign COL[13836] = 1'b0;
assign COL[13837] = 1'b0;
assign COL[13838] = 1'b0;
assign COL[13839] = 1'b0;
assign COL[13840] = 1'b0;
assign COL[13841] = 1'b0;
assign COL[13842] = 1'b0;
assign COL[13843] = 1'b0;
assign COL[13844] = 1'b0;
assign COL[13845] = 1'b0;
assign COL[13846] = 1'b0;
assign COL[13847] = 1'b0;
assign COL[13848] = 1'b0;
assign COL[13849] = 1'b0;
assign COL[13850] = 1'b1;
assign COL[13851] = 1'b1;
assign COL[13852] = 1'b1;
assign COL[13853] = 1'b1;
assign COL[13854] = 1'b1;
assign COL[13855] = 1'b0;
assign COL[13856] = 1'b0;
assign COL[13857] = 1'b0;
assign COL[13858] = 1'b0;
assign COL[13859] = 1'b0;
assign COL[13860] = 1'b0;
assign COL[13861] = 1'b0;
assign COL[13862] = 1'b0;
assign COL[13863] = 1'b0;
assign COL[13864] = 1'b0;
assign COL[13865] = 1'b0;
assign COL[13866] = 1'b0;
assign COL[13867] = 1'b0;
assign COL[13868] = 1'b0;
assign COL[13869] = 1'b0;
assign COL[13870] = 1'b0;
assign COL[13871] = 1'b0;
assign COL[13872] = 1'b0;
assign COL[13873] = 1'b0;
assign COL[13874] = 1'b0;
assign COL[13875] = 1'b0;
assign COL[13876] = 1'b0;
assign COL[13877] = 1'b0;
assign COL[13878] = 1'b0;
assign COL[13879] = 1'b0;
assign COL[13880] = 1'b0;
assign COL[13881] = 1'b0;
assign COL[13882] = 1'b0;
assign COL[13883] = 1'b0;
assign COL[13884] = 1'b0;
assign COL[13885] = 1'b0;
assign COL[13886] = 1'b0;
assign COL[13887] = 1'b0;
assign COL[13888] = 1'b0;
assign COL[13889] = 1'b0;
assign COL[13890] = 1'b0;
assign COL[13891] = 1'b0;
assign COL[13892] = 1'b0;
assign COL[13893] = 1'b0;
assign COL[13894] = 1'b0;
assign COL[13895] = 1'b0;
assign COL[13896] = 1'b0;
assign COL[13897] = 1'b0;
assign COL[13898] = 1'b0;
assign COL[13899] = 1'b0;
assign COL[13900] = 1'b0;
assign COL[13901] = 1'b0;
assign COL[13902] = 1'b0;
assign COL[13903] = 1'b0;
assign COL[13904] = 1'b0;
assign COL[13905] = 1'b0;
assign COL[13906] = 1'b0;
assign COL[13907] = 1'b0;
assign COL[13908] = 1'b0;
assign COL[13909] = 1'b0;
assign COL[13910] = 1'b0;
assign COL[13911] = 1'b0;
assign COL[13912] = 1'b0;
assign COL[13913] = 1'b0;
assign COL[13914] = 1'b0;
assign COL[13915] = 1'b0;
assign COL[13916] = 1'b0;
assign COL[13917] = 1'b0;
assign COL[13918] = 1'b0;
assign COL[13919] = 1'b0;
assign COL[13920] = 1'b0;
assign COL[13921] = 1'b1;
assign COL[13922] = 1'b1;
assign COL[13923] = 1'b1;
assign COL[13924] = 1'b1;
assign COL[13925] = 1'b0;
assign COL[13926] = 1'b0;
assign COL[13927] = 1'b0;
assign COL[13928] = 1'b0;
assign COL[13929] = 1'b0;
assign COL[13930] = 1'b0;
assign COL[13931] = 1'b0;
assign COL[13932] = 1'b0;
assign COL[13933] = 1'b0;
assign COL[13934] = 1'b0;
assign COL[13935] = 1'b0;
assign COL[13936] = 1'b0;
assign COL[13937] = 1'b0;
assign COL[13938] = 1'b0;
assign COL[13939] = 1'b0;
assign COL[13940] = 1'b0;
assign COL[13941] = 1'b0;
assign COL[13942] = 1'b0;
assign COL[13943] = 1'b0;
assign COL[13944] = 1'b0;
assign COL[13945] = 1'b0;
assign COL[13946] = 1'b0;
assign COL[13947] = 1'b0;
assign COL[13948] = 1'b0;
assign COL[13949] = 1'b0;
assign COL[13950] = 1'b0;
assign COL[13951] = 1'b0;
assign COL[13952] = 1'b0;
assign COL[13953] = 1'b0;
assign COL[13954] = 1'b0;
assign COL[13955] = 1'b0;
assign COL[13956] = 1'b0;
assign COL[13957] = 1'b0;
assign COL[13958] = 1'b0;
assign COL[13959] = 1'b0;
assign COL[13960] = 1'b0;
assign COL[13961] = 1'b0;
assign COL[13962] = 1'b0;
assign COL[13963] = 1'b0;
assign COL[13964] = 1'b0;
assign COL[13965] = 1'b0;
assign COL[13966] = 1'b0;
assign COL[13967] = 1'b0;
assign COL[13968] = 1'b0;
assign COL[13969] = 1'b0;
assign COL[13970] = 1'b0;
assign COL[13971] = 1'b0;
assign COL[13972] = 1'b0;
assign COL[13973] = 1'b0;
assign COL[13974] = 1'b0;
assign COL[13975] = 1'b1;
assign COL[13976] = 1'b1;
assign COL[13977] = 1'b1;
assign COL[13978] = 1'b1;
assign COL[13979] = 1'b0;
assign COL[13980] = 1'b0;
assign COL[13981] = 1'b0;
assign COL[13982] = 1'b0;
assign COL[13983] = 1'b0;
assign COL[13984] = 1'b0;
assign COL[13985] = 1'b0;
assign COL[13986] = 1'b0;
assign COL[13987] = 1'b0;
assign COL[13988] = 1'b0;
assign COL[13989] = 1'b0;
assign COL[13990] = 1'b0;
assign COL[13991] = 1'b0;
assign COL[13992] = 1'b0;
assign COL[13993] = 1'b0;
assign COL[13994] = 1'b0;
assign COL[13995] = 1'b0;
assign COL[13996] = 1'b0;
assign COL[13997] = 1'b0;
assign COL[13998] = 1'b0;
assign COL[13999] = 1'b0;
assign COL[14000] = 1'b0;
assign COL[14001] = 1'b0;
assign COL[14002] = 1'b0;
assign COL[14003] = 1'b0;
assign COL[14004] = 1'b0;
assign COL[14005] = 1'b0;
assign COL[14006] = 1'b0;
assign COL[14007] = 1'b0;
assign COL[14008] = 1'b0;
assign COL[14009] = 1'b0;
assign COL[14010] = 1'b1;
assign COL[14011] = 1'b1;
assign COL[14012] = 1'b1;
assign COL[14013] = 1'b1;
assign COL[14014] = 1'b1;
assign COL[14015] = 1'b0;
assign COL[14016] = 1'b0;
assign COL[14017] = 1'b0;
assign COL[14018] = 1'b0;
assign COL[14019] = 1'b0;
assign COL[14020] = 1'b0;
assign COL[14021] = 1'b0;
assign COL[14022] = 1'b0;
assign COL[14023] = 1'b0;
assign COL[14024] = 1'b0;
assign COL[14025] = 1'b0;
assign COL[14026] = 1'b0;
assign COL[14027] = 1'b0;
assign COL[14028] = 1'b0;
assign COL[14029] = 1'b0;
assign COL[14030] = 1'b0;
assign COL[14031] = 1'b0;
assign COL[14032] = 1'b0;
assign COL[14033] = 1'b0;
assign COL[14034] = 1'b0;
assign COL[14035] = 1'b0;
assign COL[14036] = 1'b0;
assign COL[14037] = 1'b0;
assign COL[14038] = 1'b0;
assign COL[14039] = 1'b0;
assign COL[14040] = 1'b0;
assign COL[14041] = 1'b0;
assign COL[14042] = 1'b0;
assign COL[14043] = 1'b0;
assign COL[14044] = 1'b0;
assign COL[14045] = 1'b0;
assign COL[14046] = 1'b0;
assign COL[14047] = 1'b0;
assign COL[14048] = 1'b0;
assign COL[14049] = 1'b0;
assign COL[14050] = 1'b0;
assign COL[14051] = 1'b0;
assign COL[14052] = 1'b0;
assign COL[14053] = 1'b0;
assign COL[14054] = 1'b0;
assign COL[14055] = 1'b0;
assign COL[14056] = 1'b0;
assign COL[14057] = 1'b0;
assign COL[14058] = 1'b0;
assign COL[14059] = 1'b0;
assign COL[14060] = 1'b0;
assign COL[14061] = 1'b0;
assign COL[14062] = 1'b0;
assign COL[14063] = 1'b0;
assign COL[14064] = 1'b0;
assign COL[14065] = 1'b0;
assign COL[14066] = 1'b0;
assign COL[14067] = 1'b0;
assign COL[14068] = 1'b0;
assign COL[14069] = 1'b0;
assign COL[14070] = 1'b0;
assign COL[14071] = 1'b0;
assign COL[14072] = 1'b0;
assign COL[14073] = 1'b0;
assign COL[14074] = 1'b0;
assign COL[14075] = 1'b0;
assign COL[14076] = 1'b0;
assign COL[14077] = 1'b0;
assign COL[14078] = 1'b0;
assign COL[14079] = 1'b0;
assign COL[14080] = 1'b0;
assign COL[14081] = 1'b1;
assign COL[14082] = 1'b1;
assign COL[14083] = 1'b1;
assign COL[14084] = 1'b1;
assign COL[14085] = 1'b0;
assign COL[14086] = 1'b0;
assign COL[14087] = 1'b0;
assign COL[14088] = 1'b0;
assign COL[14089] = 1'b0;
assign COL[14090] = 1'b0;
assign COL[14091] = 1'b0;
assign COL[14092] = 1'b0;
assign COL[14093] = 1'b0;
assign COL[14094] = 1'b0;
assign COL[14095] = 1'b0;
assign COL[14096] = 1'b0;
assign COL[14097] = 1'b0;
assign COL[14098] = 1'b0;
assign COL[14099] = 1'b0;
assign COL[14100] = 1'b0;
assign COL[14101] = 1'b0;
assign COL[14102] = 1'b0;
assign COL[14103] = 1'b0;
assign COL[14104] = 1'b0;
assign COL[14105] = 1'b0;
assign COL[14106] = 1'b0;
assign COL[14107] = 1'b0;
assign COL[14108] = 1'b0;
assign COL[14109] = 1'b0;
assign COL[14110] = 1'b0;
assign COL[14111] = 1'b0;
assign COL[14112] = 1'b0;
assign COL[14113] = 1'b0;
assign COL[14114] = 1'b0;
assign COL[14115] = 1'b0;
assign COL[14116] = 1'b0;
assign COL[14117] = 1'b0;
assign COL[14118] = 1'b0;
assign COL[14119] = 1'b0;
assign COL[14120] = 1'b0;
assign COL[14121] = 1'b0;
assign COL[14122] = 1'b0;
assign COL[14123] = 1'b0;
assign COL[14124] = 1'b0;
assign COL[14125] = 1'b0;
assign COL[14126] = 1'b0;
assign COL[14127] = 1'b0;
assign COL[14128] = 1'b0;
assign COL[14129] = 1'b0;
assign COL[14130] = 1'b0;
assign COL[14131] = 1'b0;
assign COL[14132] = 1'b0;
assign COL[14133] = 1'b0;
assign COL[14134] = 1'b0;
assign COL[14135] = 1'b1;
assign COL[14136] = 1'b1;
assign COL[14137] = 1'b1;
assign COL[14138] = 1'b1;
assign COL[14139] = 1'b0;
assign COL[14140] = 1'b0;
assign COL[14141] = 1'b0;
assign COL[14142] = 1'b0;
assign COL[14143] = 1'b0;
assign COL[14144] = 1'b0;
assign COL[14145] = 1'b0;
assign COL[14146] = 1'b0;
assign COL[14147] = 1'b0;
assign COL[14148] = 1'b0;
assign COL[14149] = 1'b0;
assign COL[14150] = 1'b0;
assign COL[14151] = 1'b0;
assign COL[14152] = 1'b0;
assign COL[14153] = 1'b0;
assign COL[14154] = 1'b0;
assign COL[14155] = 1'b0;
assign COL[14156] = 1'b0;
assign COL[14157] = 1'b0;
assign COL[14158] = 1'b0;
assign COL[14159] = 1'b0;
assign COL[14160] = 1'b0;
assign COL[14161] = 1'b0;
assign COL[14162] = 1'b0;
assign COL[14163] = 1'b0;
assign COL[14164] = 1'b0;
assign COL[14165] = 1'b0;
assign COL[14166] = 1'b0;
assign COL[14167] = 1'b0;
assign COL[14168] = 1'b0;
assign COL[14169] = 1'b0;
assign COL[14170] = 1'b1;
assign COL[14171] = 1'b1;
assign COL[14172] = 1'b1;
assign COL[14173] = 1'b1;
assign COL[14174] = 1'b1;
assign COL[14175] = 1'b0;
assign COL[14176] = 1'b0;
assign COL[14177] = 1'b0;
assign COL[14178] = 1'b0;
assign COL[14179] = 1'b0;
assign COL[14180] = 1'b0;
assign COL[14181] = 1'b0;
assign COL[14182] = 1'b0;
assign COL[14183] = 1'b0;
assign COL[14184] = 1'b0;
assign COL[14185] = 1'b0;
assign COL[14186] = 1'b0;
assign COL[14187] = 1'b0;
assign COL[14188] = 1'b0;
assign COL[14189] = 1'b0;
assign COL[14190] = 1'b0;
assign COL[14191] = 1'b0;
assign COL[14192] = 1'b0;
assign COL[14193] = 1'b0;
assign COL[14194] = 1'b0;
assign COL[14195] = 1'b0;
assign COL[14196] = 1'b0;
assign COL[14197] = 1'b0;
assign COL[14198] = 1'b0;
assign COL[14199] = 1'b0;
assign COL[14200] = 1'b0;
assign COL[14201] = 1'b0;
assign COL[14202] = 1'b0;
assign COL[14203] = 1'b0;
assign COL[14204] = 1'b0;
assign COL[14205] = 1'b0;
assign COL[14206] = 1'b0;
assign COL[14207] = 1'b0;
assign COL[14208] = 1'b0;
assign COL[14209] = 1'b0;
assign COL[14210] = 1'b0;
assign COL[14211] = 1'b0;
assign COL[14212] = 1'b0;
assign COL[14213] = 1'b0;
assign COL[14214] = 1'b0;
assign COL[14215] = 1'b0;
assign COL[14216] = 1'b0;
assign COL[14217] = 1'b0;
assign COL[14218] = 1'b0;
assign COL[14219] = 1'b0;
assign COL[14220] = 1'b0;
assign COL[14221] = 1'b0;
assign COL[14222] = 1'b0;
assign COL[14223] = 1'b0;
assign COL[14224] = 1'b0;
assign COL[14225] = 1'b0;
assign COL[14226] = 1'b0;
assign COL[14227] = 1'b0;
assign COL[14228] = 1'b0;
assign COL[14229] = 1'b0;
assign COL[14230] = 1'b0;
assign COL[14231] = 1'b0;
assign COL[14232] = 1'b0;
assign COL[14233] = 1'b0;
assign COL[14234] = 1'b0;
assign COL[14235] = 1'b0;
assign COL[14236] = 1'b0;
assign COL[14237] = 1'b0;
assign COL[14238] = 1'b0;
assign COL[14239] = 1'b0;
assign COL[14240] = 1'b0;
assign COL[14241] = 1'b1;
assign COL[14242] = 1'b1;
assign COL[14243] = 1'b1;
assign COL[14244] = 1'b1;
assign COL[14245] = 1'b1;
assign COL[14246] = 1'b1;
assign COL[14247] = 1'b1;
assign COL[14248] = 1'b1;
assign COL[14249] = 1'b1;
assign COL[14250] = 1'b1;
assign COL[14251] = 1'b1;
assign COL[14252] = 1'b1;
assign COL[14253] = 1'b1;
assign COL[14254] = 1'b1;
assign COL[14255] = 1'b1;
assign COL[14256] = 1'b1;
assign COL[14257] = 1'b1;
assign COL[14258] = 1'b1;
assign COL[14259] = 1'b1;
assign COL[14260] = 1'b1;
assign COL[14261] = 1'b1;
assign COL[14262] = 1'b1;
assign COL[14263] = 1'b1;
assign COL[14264] = 1'b1;
assign COL[14265] = 1'b1;
assign COL[14266] = 1'b1;
assign COL[14267] = 1'b1;
assign COL[14268] = 1'b1;
assign COL[14269] = 1'b1;
assign COL[14270] = 1'b1;
assign COL[14271] = 1'b1;
assign COL[14272] = 1'b1;
assign COL[14273] = 1'b1;
assign COL[14274] = 1'b1;
assign COL[14275] = 1'b1;
assign COL[14276] = 1'b1;
assign COL[14277] = 1'b1;
assign COL[14278] = 1'b1;
assign COL[14279] = 1'b1;
assign COL[14280] = 1'b1;
assign COL[14281] = 1'b1;
assign COL[14282] = 1'b1;
assign COL[14283] = 1'b1;
assign COL[14284] = 1'b1;
assign COL[14285] = 1'b1;
assign COL[14286] = 1'b1;
assign COL[14287] = 1'b1;
assign COL[14288] = 1'b1;
assign COL[14289] = 1'b1;
assign COL[14290] = 1'b1;
assign COL[14291] = 1'b1;
assign COL[14292] = 1'b1;
assign COL[14293] = 1'b1;
assign COL[14294] = 1'b1;
assign COL[14295] = 1'b1;
assign COL[14296] = 1'b1;
assign COL[14297] = 1'b1;
assign COL[14298] = 1'b1;
assign COL[14299] = 1'b1;
assign COL[14300] = 1'b1;
assign COL[14301] = 1'b1;
assign COL[14302] = 1'b1;
assign COL[14303] = 1'b1;
assign COL[14304] = 1'b1;
assign COL[14305] = 1'b1;
assign COL[14306] = 1'b1;
assign COL[14307] = 1'b1;
assign COL[14308] = 1'b1;
assign COL[14309] = 1'b1;
assign COL[14310] = 1'b1;
assign COL[14311] = 1'b1;
assign COL[14312] = 1'b1;
assign COL[14313] = 1'b1;
assign COL[14314] = 1'b1;
assign COL[14315] = 1'b1;
assign COL[14316] = 1'b1;
assign COL[14317] = 1'b1;
assign COL[14318] = 1'b1;
assign COL[14319] = 1'b1;
assign COL[14320] = 1'b1;
assign COL[14321] = 1'b1;
assign COL[14322] = 1'b1;
assign COL[14323] = 1'b1;
assign COL[14324] = 1'b1;
assign COL[14325] = 1'b1;
assign COL[14326] = 1'b1;
assign COL[14327] = 1'b1;
assign COL[14328] = 1'b1;
assign COL[14329] = 1'b1;
assign COL[14330] = 1'b1;
assign COL[14331] = 1'b1;
assign COL[14332] = 1'b1;
assign COL[14333] = 1'b1;
assign COL[14334] = 1'b1;
assign COL[14335] = 1'b0;
assign COL[14336] = 1'b0;
assign COL[14337] = 1'b0;
assign COL[14338] = 1'b0;
assign COL[14339] = 1'b0;
assign COL[14340] = 1'b0;
assign COL[14341] = 1'b0;
assign COL[14342] = 1'b0;
assign COL[14343] = 1'b0;
assign COL[14344] = 1'b0;
assign COL[14345] = 1'b0;
assign COL[14346] = 1'b0;
assign COL[14347] = 1'b0;
assign COL[14348] = 1'b0;
assign COL[14349] = 1'b0;
assign COL[14350] = 1'b0;
assign COL[14351] = 1'b0;
assign COL[14352] = 1'b0;
assign COL[14353] = 1'b0;
assign COL[14354] = 1'b0;
assign COL[14355] = 1'b0;
assign COL[14356] = 1'b0;
assign COL[14357] = 1'b0;
assign COL[14358] = 1'b0;
assign COL[14359] = 1'b0;
assign COL[14360] = 1'b0;
assign COL[14361] = 1'b0;
assign COL[14362] = 1'b0;
assign COL[14363] = 1'b0;
assign COL[14364] = 1'b0;
assign COL[14365] = 1'b0;
assign COL[14366] = 1'b0;
assign COL[14367] = 1'b0;
assign COL[14368] = 1'b0;
assign COL[14369] = 1'b0;
assign COL[14370] = 1'b0;
assign COL[14371] = 1'b0;
assign COL[14372] = 1'b0;
assign COL[14373] = 1'b0;
assign COL[14374] = 1'b0;
assign COL[14375] = 1'b0;
assign COL[14376] = 1'b0;
assign COL[14377] = 1'b0;
assign COL[14378] = 1'b0;
assign COL[14379] = 1'b0;
assign COL[14380] = 1'b0;
assign COL[14381] = 1'b0;
assign COL[14382] = 1'b0;
assign COL[14383] = 1'b0;
assign COL[14384] = 1'b0;
assign COL[14385] = 1'b0;
assign COL[14386] = 1'b0;
assign COL[14387] = 1'b0;
assign COL[14388] = 1'b0;
assign COL[14389] = 1'b0;
assign COL[14390] = 1'b0;
assign COL[14391] = 1'b0;
assign COL[14392] = 1'b0;
assign COL[14393] = 1'b0;
assign COL[14394] = 1'b0;
assign COL[14395] = 1'b0;
assign COL[14396] = 1'b0;
assign COL[14397] = 1'b0;
assign COL[14398] = 1'b0;
assign COL[14399] = 1'b0;
assign COL[14400] = 1'b0;
assign COL[14401] = 1'b1;
assign COL[14402] = 1'b1;
assign COL[14403] = 1'b1;
assign COL[14404] = 1'b1;
assign COL[14405] = 1'b1;
assign COL[14406] = 1'b1;
assign COL[14407] = 1'b1;
assign COL[14408] = 1'b1;
assign COL[14409] = 1'b1;
assign COL[14410] = 1'b1;
assign COL[14411] = 1'b1;
assign COL[14412] = 1'b1;
assign COL[14413] = 1'b1;
assign COL[14414] = 1'b1;
assign COL[14415] = 1'b1;
assign COL[14416] = 1'b1;
assign COL[14417] = 1'b1;
assign COL[14418] = 1'b1;
assign COL[14419] = 1'b1;
assign COL[14420] = 1'b1;
assign COL[14421] = 1'b1;
assign COL[14422] = 1'b1;
assign COL[14423] = 1'b1;
assign COL[14424] = 1'b1;
assign COL[14425] = 1'b1;
assign COL[14426] = 1'b1;
assign COL[14427] = 1'b1;
assign COL[14428] = 1'b1;
assign COL[14429] = 1'b1;
assign COL[14430] = 1'b1;
assign COL[14431] = 1'b1;
assign COL[14432] = 1'b1;
assign COL[14433] = 1'b1;
assign COL[14434] = 1'b1;
assign COL[14435] = 1'b1;
assign COL[14436] = 1'b1;
assign COL[14437] = 1'b1;
assign COL[14438] = 1'b1;
assign COL[14439] = 1'b1;
assign COL[14440] = 1'b1;
assign COL[14441] = 1'b1;
assign COL[14442] = 1'b1;
assign COL[14443] = 1'b1;
assign COL[14444] = 1'b1;
assign COL[14445] = 1'b1;
assign COL[14446] = 1'b1;
assign COL[14447] = 1'b1;
assign COL[14448] = 1'b1;
assign COL[14449] = 1'b1;
assign COL[14450] = 1'b1;
assign COL[14451] = 1'b1;
assign COL[14452] = 1'b1;
assign COL[14453] = 1'b1;
assign COL[14454] = 1'b1;
assign COL[14455] = 1'b1;
assign COL[14456] = 1'b1;
assign COL[14457] = 1'b1;
assign COL[14458] = 1'b1;
assign COL[14459] = 1'b1;
assign COL[14460] = 1'b1;
assign COL[14461] = 1'b1;
assign COL[14462] = 1'b1;
assign COL[14463] = 1'b1;
assign COL[14464] = 1'b1;
assign COL[14465] = 1'b1;
assign COL[14466] = 1'b1;
assign COL[14467] = 1'b1;
assign COL[14468] = 1'b1;
assign COL[14469] = 1'b1;
assign COL[14470] = 1'b1;
assign COL[14471] = 1'b1;
assign COL[14472] = 1'b1;
assign COL[14473] = 1'b1;
assign COL[14474] = 1'b1;
assign COL[14475] = 1'b1;
assign COL[14476] = 1'b1;
assign COL[14477] = 1'b1;
assign COL[14478] = 1'b1;
assign COL[14479] = 1'b1;
assign COL[14480] = 1'b1;
assign COL[14481] = 1'b1;
assign COL[14482] = 1'b1;
assign COL[14483] = 1'b1;
assign COL[14484] = 1'b1;
assign COL[14485] = 1'b1;
assign COL[14486] = 1'b1;
assign COL[14487] = 1'b1;
assign COL[14488] = 1'b1;
assign COL[14489] = 1'b1;
assign COL[14490] = 1'b1;
assign COL[14491] = 1'b1;
assign COL[14492] = 1'b1;
assign COL[14493] = 1'b1;
assign COL[14494] = 1'b1;
assign COL[14495] = 1'b0;
assign COL[14496] = 1'b0;
assign COL[14497] = 1'b0;
assign COL[14498] = 1'b0;
assign COL[14499] = 1'b0;
assign COL[14500] = 1'b0;
assign COL[14501] = 1'b0;
assign COL[14502] = 1'b0;
assign COL[14503] = 1'b0;
assign COL[14504] = 1'b0;
assign COL[14505] = 1'b0;
assign COL[14506] = 1'b0;
assign COL[14507] = 1'b0;
assign COL[14508] = 1'b0;
assign COL[14509] = 1'b0;
assign COL[14510] = 1'b0;
assign COL[14511] = 1'b0;
assign COL[14512] = 1'b0;
assign COL[14513] = 1'b0;
assign COL[14514] = 1'b0;
assign COL[14515] = 1'b0;
assign COL[14516] = 1'b0;
assign COL[14517] = 1'b0;
assign COL[14518] = 1'b0;
assign COL[14519] = 1'b0;
assign COL[14520] = 1'b0;
assign COL[14521] = 1'b0;
assign COL[14522] = 1'b0;
assign COL[14523] = 1'b0;
assign COL[14524] = 1'b0;
assign COL[14525] = 1'b0;
assign COL[14526] = 1'b0;
assign COL[14527] = 1'b0;
assign COL[14528] = 1'b0;
assign COL[14529] = 1'b0;
assign COL[14530] = 1'b0;
assign COL[14531] = 1'b0;
assign COL[14532] = 1'b0;
assign COL[14533] = 1'b0;
assign COL[14534] = 1'b0;
assign COL[14535] = 1'b0;
assign COL[14536] = 1'b0;
assign COL[14537] = 1'b0;
assign COL[14538] = 1'b0;
assign COL[14539] = 1'b0;
assign COL[14540] = 1'b0;
assign COL[14541] = 1'b0;
assign COL[14542] = 1'b0;
assign COL[14543] = 1'b0;
assign COL[14544] = 1'b0;
assign COL[14545] = 1'b0;
assign COL[14546] = 1'b0;
assign COL[14547] = 1'b0;
assign COL[14548] = 1'b0;
assign COL[14549] = 1'b0;
assign COL[14550] = 1'b0;
assign COL[14551] = 1'b0;
assign COL[14552] = 1'b0;
assign COL[14553] = 1'b0;
assign COL[14554] = 1'b0;
assign COL[14555] = 1'b0;
assign COL[14556] = 1'b0;
assign COL[14557] = 1'b0;
assign COL[14558] = 1'b0;
assign COL[14559] = 1'b0;
assign COL[14560] = 1'b0;
assign COL[14561] = 1'b1;
assign COL[14562] = 1'b1;
assign COL[14563] = 1'b1;
assign COL[14564] = 1'b1;
assign COL[14565] = 1'b1;
assign COL[14566] = 1'b1;
assign COL[14567] = 1'b1;
assign COL[14568] = 1'b1;
assign COL[14569] = 1'b1;
assign COL[14570] = 1'b1;
assign COL[14571] = 1'b1;
assign COL[14572] = 1'b1;
assign COL[14573] = 1'b1;
assign COL[14574] = 1'b1;
assign COL[14575] = 1'b1;
assign COL[14576] = 1'b1;
assign COL[14577] = 1'b1;
assign COL[14578] = 1'b1;
assign COL[14579] = 1'b1;
assign COL[14580] = 1'b1;
assign COL[14581] = 1'b1;
assign COL[14582] = 1'b1;
assign COL[14583] = 1'b1;
assign COL[14584] = 1'b1;
assign COL[14585] = 1'b1;
assign COL[14586] = 1'b1;
assign COL[14587] = 1'b1;
assign COL[14588] = 1'b1;
assign COL[14589] = 1'b1;
assign COL[14590] = 1'b1;
assign COL[14591] = 1'b1;
assign COL[14592] = 1'b1;
assign COL[14593] = 1'b1;
assign COL[14594] = 1'b1;
assign COL[14595] = 1'b1;
assign COL[14596] = 1'b1;
assign COL[14597] = 1'b1;
assign COL[14598] = 1'b1;
assign COL[14599] = 1'b1;
assign COL[14600] = 1'b1;
assign COL[14601] = 1'b1;
assign COL[14602] = 1'b1;
assign COL[14603] = 1'b1;
assign COL[14604] = 1'b1;
assign COL[14605] = 1'b1;
assign COL[14606] = 1'b1;
assign COL[14607] = 1'b1;
assign COL[14608] = 1'b1;
assign COL[14609] = 1'b1;
assign COL[14610] = 1'b1;
assign COL[14611] = 1'b1;
assign COL[14612] = 1'b1;
assign COL[14613] = 1'b1;
assign COL[14614] = 1'b1;
assign COL[14615] = 1'b1;
assign COL[14616] = 1'b1;
assign COL[14617] = 1'b1;
assign COL[14618] = 1'b1;
assign COL[14619] = 1'b1;
assign COL[14620] = 1'b1;
assign COL[14621] = 1'b1;
assign COL[14622] = 1'b1;
assign COL[14623] = 1'b1;
assign COL[14624] = 1'b1;
assign COL[14625] = 1'b1;
assign COL[14626] = 1'b1;
assign COL[14627] = 1'b1;
assign COL[14628] = 1'b1;
assign COL[14629] = 1'b1;
assign COL[14630] = 1'b1;
assign COL[14631] = 1'b1;
assign COL[14632] = 1'b1;
assign COL[14633] = 1'b1;
assign COL[14634] = 1'b1;
assign COL[14635] = 1'b1;
assign COL[14636] = 1'b1;
assign COL[14637] = 1'b1;
assign COL[14638] = 1'b1;
assign COL[14639] = 1'b1;
assign COL[14640] = 1'b1;
assign COL[14641] = 1'b1;
assign COL[14642] = 1'b1;
assign COL[14643] = 1'b1;
assign COL[14644] = 1'b1;
assign COL[14645] = 1'b1;
assign COL[14646] = 1'b1;
assign COL[14647] = 1'b1;
assign COL[14648] = 1'b1;
assign COL[14649] = 1'b1;
assign COL[14650] = 1'b1;
assign COL[14651] = 1'b1;
assign COL[14652] = 1'b1;
assign COL[14653] = 1'b1;
assign COL[14654] = 1'b1;
assign COL[14655] = 1'b0;
assign COL[14656] = 1'b0;
assign COL[14657] = 1'b0;
assign COL[14658] = 1'b0;
assign COL[14659] = 1'b0;
assign COL[14660] = 1'b0;
assign COL[14661] = 1'b0;
assign COL[14662] = 1'b0;
assign COL[14663] = 1'b0;
assign COL[14664] = 1'b0;
assign COL[14665] = 1'b0;
assign COL[14666] = 1'b0;
assign COL[14667] = 1'b0;
assign COL[14668] = 1'b0;
assign COL[14669] = 1'b0;
assign COL[14670] = 1'b0;
assign COL[14671] = 1'b0;
assign COL[14672] = 1'b0;
assign COL[14673] = 1'b0;
assign COL[14674] = 1'b0;
assign COL[14675] = 1'b0;
assign COL[14676] = 1'b0;
assign COL[14677] = 1'b0;
assign COL[14678] = 1'b0;
assign COL[14679] = 1'b0;
assign COL[14680] = 1'b0;
assign COL[14681] = 1'b0;
assign COL[14682] = 1'b0;
assign COL[14683] = 1'b0;
assign COL[14684] = 1'b0;
assign COL[14685] = 1'b0;
assign COL[14686] = 1'b0;
assign COL[14687] = 1'b0;
assign COL[14688] = 1'b0;
assign COL[14689] = 1'b0;
assign COL[14690] = 1'b0;
assign COL[14691] = 1'b0;
assign COL[14692] = 1'b0;
assign COL[14693] = 1'b0;
assign COL[14694] = 1'b0;
assign COL[14695] = 1'b0;
assign COL[14696] = 1'b0;
assign COL[14697] = 1'b0;
assign COL[14698] = 1'b0;
assign COL[14699] = 1'b0;
assign COL[14700] = 1'b0;
assign COL[14701] = 1'b0;
assign COL[14702] = 1'b0;
assign COL[14703] = 1'b0;
assign COL[14704] = 1'b0;
assign COL[14705] = 1'b0;
assign COL[14706] = 1'b0;
assign COL[14707] = 1'b0;
assign COL[14708] = 1'b0;
assign COL[14709] = 1'b0;
assign COL[14710] = 1'b0;
assign COL[14711] = 1'b0;
assign COL[14712] = 1'b0;
assign COL[14713] = 1'b0;
assign COL[14714] = 1'b0;
assign COL[14715] = 1'b0;
assign COL[14716] = 1'b0;
assign COL[14717] = 1'b0;
assign COL[14718] = 1'b0;
assign COL[14719] = 1'b0;
assign COL[14720] = 1'b0;
assign COL[14721] = 1'b1;
assign COL[14722] = 1'b1;
assign COL[14723] = 1'b1;
assign COL[14724] = 1'b1;
assign COL[14725] = 1'b1;
assign COL[14726] = 1'b1;
assign COL[14727] = 1'b1;
assign COL[14728] = 1'b1;
assign COL[14729] = 1'b1;
assign COL[14730] = 1'b1;
assign COL[14731] = 1'b1;
assign COL[14732] = 1'b1;
assign COL[14733] = 1'b1;
assign COL[14734] = 1'b1;
assign COL[14735] = 1'b1;
assign COL[14736] = 1'b1;
assign COL[14737] = 1'b1;
assign COL[14738] = 1'b1;
assign COL[14739] = 1'b1;
assign COL[14740] = 1'b1;
assign COL[14741] = 1'b1;
assign COL[14742] = 1'b1;
assign COL[14743] = 1'b1;
assign COL[14744] = 1'b1;
assign COL[14745] = 1'b1;
assign COL[14746] = 1'b1;
assign COL[14747] = 1'b1;
assign COL[14748] = 1'b1;
assign COL[14749] = 1'b1;
assign COL[14750] = 1'b1;
assign COL[14751] = 1'b1;
assign COL[14752] = 1'b1;
assign COL[14753] = 1'b1;
assign COL[14754] = 1'b1;
assign COL[14755] = 1'b1;
assign COL[14756] = 1'b1;
assign COL[14757] = 1'b1;
assign COL[14758] = 1'b1;
assign COL[14759] = 1'b1;
assign COL[14760] = 1'b1;
assign COL[14761] = 1'b1;
assign COL[14762] = 1'b1;
assign COL[14763] = 1'b1;
assign COL[14764] = 1'b1;
assign COL[14765] = 1'b1;
assign COL[14766] = 1'b1;
assign COL[14767] = 1'b1;
assign COL[14768] = 1'b1;
assign COL[14769] = 1'b1;
assign COL[14770] = 1'b1;
assign COL[14771] = 1'b1;
assign COL[14772] = 1'b1;
assign COL[14773] = 1'b1;
assign COL[14774] = 1'b1;
assign COL[14775] = 1'b1;
assign COL[14776] = 1'b1;
assign COL[14777] = 1'b1;
assign COL[14778] = 1'b1;
assign COL[14779] = 1'b1;
assign COL[14780] = 1'b1;
assign COL[14781] = 1'b1;
assign COL[14782] = 1'b1;
assign COL[14783] = 1'b1;
assign COL[14784] = 1'b1;
assign COL[14785] = 1'b1;
assign COL[14786] = 1'b1;
assign COL[14787] = 1'b1;
assign COL[14788] = 1'b1;
assign COL[14789] = 1'b1;
assign COL[14790] = 1'b1;
assign COL[14791] = 1'b1;
assign COL[14792] = 1'b1;
assign COL[14793] = 1'b1;
assign COL[14794] = 1'b1;
assign COL[14795] = 1'b1;
assign COL[14796] = 1'b1;
assign COL[14797] = 1'b1;
assign COL[14798] = 1'b1;
assign COL[14799] = 1'b1;
assign COL[14800] = 1'b1;
assign COL[14801] = 1'b1;
assign COL[14802] = 1'b1;
assign COL[14803] = 1'b1;
assign COL[14804] = 1'b1;
assign COL[14805] = 1'b1;
assign COL[14806] = 1'b1;
assign COL[14807] = 1'b1;
assign COL[14808] = 1'b1;
assign COL[14809] = 1'b1;
assign COL[14810] = 1'b1;
assign COL[14811] = 1'b1;
assign COL[14812] = 1'b1;
assign COL[14813] = 1'b1;
assign COL[14814] = 1'b1;
assign COL[14815] = 1'b0;
assign COL[14816] = 1'b0;
assign COL[14817] = 1'b0;
assign COL[14818] = 1'b0;
assign COL[14819] = 1'b0;
assign COL[14820] = 1'b0;
assign COL[14821] = 1'b0;
assign COL[14822] = 1'b0;
assign COL[14823] = 1'b0;
assign COL[14824] = 1'b0;
assign COL[14825] = 1'b0;
assign COL[14826] = 1'b0;
assign COL[14827] = 1'b0;
assign COL[14828] = 1'b0;
assign COL[14829] = 1'b0;
assign COL[14830] = 1'b0;
assign COL[14831] = 1'b0;
assign COL[14832] = 1'b0;
assign COL[14833] = 1'b0;
assign COL[14834] = 1'b0;
assign COL[14835] = 1'b0;
assign COL[14836] = 1'b0;
assign COL[14837] = 1'b0;
assign COL[14838] = 1'b0;
assign COL[14839] = 1'b0;
assign COL[14840] = 1'b0;
assign COL[14841] = 1'b0;
assign COL[14842] = 1'b0;
assign COL[14843] = 1'b0;
assign COL[14844] = 1'b0;
assign COL[14845] = 1'b0;
assign COL[14846] = 1'b0;
assign COL[14847] = 1'b0;
assign COL[14848] = 1'b0;
assign COL[14849] = 1'b0;
assign COL[14850] = 1'b0;
assign COL[14851] = 1'b0;
assign COL[14852] = 1'b0;
assign COL[14853] = 1'b0;
assign COL[14854] = 1'b0;
assign COL[14855] = 1'b0;
assign COL[14856] = 1'b0;
assign COL[14857] = 1'b0;
assign COL[14858] = 1'b0;
assign COL[14859] = 1'b0;
assign COL[14860] = 1'b0;
assign COL[14861] = 1'b0;
assign COL[14862] = 1'b0;
assign COL[14863] = 1'b0;
assign COL[14864] = 1'b0;
assign COL[14865] = 1'b0;
assign COL[14866] = 1'b0;
assign COL[14867] = 1'b0;
assign COL[14868] = 1'b0;
assign COL[14869] = 1'b0;
assign COL[14870] = 1'b0;
assign COL[14871] = 1'b0;
assign COL[14872] = 1'b0;
assign COL[14873] = 1'b0;
assign COL[14874] = 1'b0;
assign COL[14875] = 1'b0;
assign COL[14876] = 1'b0;
assign COL[14877] = 1'b0;
assign COL[14878] = 1'b0;
assign COL[14879] = 1'b0;
assign COL[14880] = 1'b0;
assign COL[14881] = 1'b0;
assign COL[14882] = 1'b0;
assign COL[14883] = 1'b0;
assign COL[14884] = 1'b0;
assign COL[14885] = 1'b0;
assign COL[14886] = 1'b0;
assign COL[14887] = 1'b0;
assign COL[14888] = 1'b0;
assign COL[14889] = 1'b0;
assign COL[14890] = 1'b0;
assign COL[14891] = 1'b0;
assign COL[14892] = 1'b0;
assign COL[14893] = 1'b0;
assign COL[14894] = 1'b0;
assign COL[14895] = 1'b0;
assign COL[14896] = 1'b0;
assign COL[14897] = 1'b0;
assign COL[14898] = 1'b0;
assign COL[14899] = 1'b0;
assign COL[14900] = 1'b0;
assign COL[14901] = 1'b0;
assign COL[14902] = 1'b0;
assign COL[14903] = 1'b0;
assign COL[14904] = 1'b0;
assign COL[14905] = 1'b0;
assign COL[14906] = 1'b0;
assign COL[14907] = 1'b0;
assign COL[14908] = 1'b0;
assign COL[14909] = 1'b0;
assign COL[14910] = 1'b0;
assign COL[14911] = 1'b0;
assign COL[14912] = 1'b0;
assign COL[14913] = 1'b0;
assign COL[14914] = 1'b0;
assign COL[14915] = 1'b0;
assign COL[14916] = 1'b0;
assign COL[14917] = 1'b0;
assign COL[14918] = 1'b0;
assign COL[14919] = 1'b0;
assign COL[14920] = 1'b0;
assign COL[14921] = 1'b0;
assign COL[14922] = 1'b0;
assign COL[14923] = 1'b0;
assign COL[14924] = 1'b0;
assign COL[14925] = 1'b0;
assign COL[14926] = 1'b0;
assign COL[14927] = 1'b0;
assign COL[14928] = 1'b0;
assign COL[14929] = 1'b0;
assign COL[14930] = 1'b0;
assign COL[14931] = 1'b0;
assign COL[14932] = 1'b0;
assign COL[14933] = 1'b0;
assign COL[14934] = 1'b0;
assign COL[14935] = 1'b0;
assign COL[14936] = 1'b0;
assign COL[14937] = 1'b0;
assign COL[14938] = 1'b0;
assign COL[14939] = 1'b0;
assign COL[14940] = 1'b0;
assign COL[14941] = 1'b0;
assign COL[14942] = 1'b0;
assign COL[14943] = 1'b0;
assign COL[14944] = 1'b0;
assign COL[14945] = 1'b0;
assign COL[14946] = 1'b0;
assign COL[14947] = 1'b0;
assign COL[14948] = 1'b0;
assign COL[14949] = 1'b0;
assign COL[14950] = 1'b0;
assign COL[14951] = 1'b0;
assign COL[14952] = 1'b0;
assign COL[14953] = 1'b0;
assign COL[14954] = 1'b0;
assign COL[14955] = 1'b0;
assign COL[14956] = 1'b0;
assign COL[14957] = 1'b0;
assign COL[14958] = 1'b0;
assign COL[14959] = 1'b0;
assign COL[14960] = 1'b0;
assign COL[14961] = 1'b0;
assign COL[14962] = 1'b0;
assign COL[14963] = 1'b0;
assign COL[14964] = 1'b0;
assign COL[14965] = 1'b0;
assign COL[14966] = 1'b0;
assign COL[14967] = 1'b0;
assign COL[14968] = 1'b0;
assign COL[14969] = 1'b0;
assign COL[14970] = 1'b0;
assign COL[14971] = 1'b0;
assign COL[14972] = 1'b0;
assign COL[14973] = 1'b0;
assign COL[14974] = 1'b0;
assign COL[14975] = 1'b0;
assign COL[14976] = 1'b0;
assign COL[14977] = 1'b0;
assign COL[14978] = 1'b0;
assign COL[14979] = 1'b0;
assign COL[14980] = 1'b0;
assign COL[14981] = 1'b0;
assign COL[14982] = 1'b0;
assign COL[14983] = 1'b0;
assign COL[14984] = 1'b0;
assign COL[14985] = 1'b0;
assign COL[14986] = 1'b0;
assign COL[14987] = 1'b0;
assign COL[14988] = 1'b0;
assign COL[14989] = 1'b0;
assign COL[14990] = 1'b0;
assign COL[14991] = 1'b0;
assign COL[14992] = 1'b0;
assign COL[14993] = 1'b0;
assign COL[14994] = 1'b0;
assign COL[14995] = 1'b0;
assign COL[14996] = 1'b0;
assign COL[14997] = 1'b0;
assign COL[14998] = 1'b0;
assign COL[14999] = 1'b0;
assign COL[15000] = 1'b0;
assign COL[15001] = 1'b0;
assign COL[15002] = 1'b0;
assign COL[15003] = 1'b0;
assign COL[15004] = 1'b0;
assign COL[15005] = 1'b0;
assign COL[15006] = 1'b0;
assign COL[15007] = 1'b0;
assign COL[15008] = 1'b0;
assign COL[15009] = 1'b0;
assign COL[15010] = 1'b0;
assign COL[15011] = 1'b0;
assign COL[15012] = 1'b0;
assign COL[15013] = 1'b0;
assign COL[15014] = 1'b0;
assign COL[15015] = 1'b0;
assign COL[15016] = 1'b0;
assign COL[15017] = 1'b0;
assign COL[15018] = 1'b0;
assign COL[15019] = 1'b0;
assign COL[15020] = 1'b0;
assign COL[15021] = 1'b0;
assign COL[15022] = 1'b0;
assign COL[15023] = 1'b0;
assign COL[15024] = 1'b0;
assign COL[15025] = 1'b0;
assign COL[15026] = 1'b0;
assign COL[15027] = 1'b0;
assign COL[15028] = 1'b0;
assign COL[15029] = 1'b0;
assign COL[15030] = 1'b0;
assign COL[15031] = 1'b0;
assign COL[15032] = 1'b0;
assign COL[15033] = 1'b0;
assign COL[15034] = 1'b0;
assign COL[15035] = 1'b0;
assign COL[15036] = 1'b0;
assign COL[15037] = 1'b0;
assign COL[15038] = 1'b0;
assign COL[15039] = 1'b0;
assign COL[15040] = 1'b0;
assign COL[15041] = 1'b0;
assign COL[15042] = 1'b0;
assign COL[15043] = 1'b0;
assign COL[15044] = 1'b0;
assign COL[15045] = 1'b0;
assign COL[15046] = 1'b0;
assign COL[15047] = 1'b0;
assign COL[15048] = 1'b0;
assign COL[15049] = 1'b0;
assign COL[15050] = 1'b0;
assign COL[15051] = 1'b0;
assign COL[15052] = 1'b0;
assign COL[15053] = 1'b0;
assign COL[15054] = 1'b0;
assign COL[15055] = 1'b0;
assign COL[15056] = 1'b0;
assign COL[15057] = 1'b0;
assign COL[15058] = 1'b0;
assign COL[15059] = 1'b0;
assign COL[15060] = 1'b0;
assign COL[15061] = 1'b0;
assign COL[15062] = 1'b0;
assign COL[15063] = 1'b0;
assign COL[15064] = 1'b0;
assign COL[15065] = 1'b0;
assign COL[15066] = 1'b0;
assign COL[15067] = 1'b0;
assign COL[15068] = 1'b0;
assign COL[15069] = 1'b0;
assign COL[15070] = 1'b0;
assign COL[15071] = 1'b0;
assign COL[15072] = 1'b0;
assign COL[15073] = 1'b0;
assign COL[15074] = 1'b0;
assign COL[15075] = 1'b0;
assign COL[15076] = 1'b0;
assign COL[15077] = 1'b0;
assign COL[15078] = 1'b0;
assign COL[15079] = 1'b0;
assign COL[15080] = 1'b0;
assign COL[15081] = 1'b0;
assign COL[15082] = 1'b0;
assign COL[15083] = 1'b0;
assign COL[15084] = 1'b0;
assign COL[15085] = 1'b0;
assign COL[15086] = 1'b0;
assign COL[15087] = 1'b0;
assign COL[15088] = 1'b0;
assign COL[15089] = 1'b0;
assign COL[15090] = 1'b0;
assign COL[15091] = 1'b0;
assign COL[15092] = 1'b0;
assign COL[15093] = 1'b0;
assign COL[15094] = 1'b0;
assign COL[15095] = 1'b0;
assign COL[15096] = 1'b0;
assign COL[15097] = 1'b0;
assign COL[15098] = 1'b0;
assign COL[15099] = 1'b0;
assign COL[15100] = 1'b0;
assign COL[15101] = 1'b0;
assign COL[15102] = 1'b0;
assign COL[15103] = 1'b0;
assign COL[15104] = 1'b0;
assign COL[15105] = 1'b0;
assign COL[15106] = 1'b0;
assign COL[15107] = 1'b0;
assign COL[15108] = 1'b0;
assign COL[15109] = 1'b0;
assign COL[15110] = 1'b0;
assign COL[15111] = 1'b0;
assign COL[15112] = 1'b0;
assign COL[15113] = 1'b0;
assign COL[15114] = 1'b0;
assign COL[15115] = 1'b0;
assign COL[15116] = 1'b0;
assign COL[15117] = 1'b0;
assign COL[15118] = 1'b0;
assign COL[15119] = 1'b0;
assign COL[15120] = 1'b0;
assign COL[15121] = 1'b0;
assign COL[15122] = 1'b0;
assign COL[15123] = 1'b0;
assign COL[15124] = 1'b0;
assign COL[15125] = 1'b0;
assign COL[15126] = 1'b0;
assign COL[15127] = 1'b0;
assign COL[15128] = 1'b0;
assign COL[15129] = 1'b0;
assign COL[15130] = 1'b0;
assign COL[15131] = 1'b0;
assign COL[15132] = 1'b0;
assign COL[15133] = 1'b0;
assign COL[15134] = 1'b0;
assign COL[15135] = 1'b0;
assign COL[15136] = 1'b0;
assign COL[15137] = 1'b0;
assign COL[15138] = 1'b0;
assign COL[15139] = 1'b0;
assign COL[15140] = 1'b0;
assign COL[15141] = 1'b0;
assign COL[15142] = 1'b0;
assign COL[15143] = 1'b0;
assign COL[15144] = 1'b0;
assign COL[15145] = 1'b0;
assign COL[15146] = 1'b0;
assign COL[15147] = 1'b0;
assign COL[15148] = 1'b0;
assign COL[15149] = 1'b0;
assign COL[15150] = 1'b0;
assign COL[15151] = 1'b0;
assign COL[15152] = 1'b0;
assign COL[15153] = 1'b0;
assign COL[15154] = 1'b0;
assign COL[15155] = 1'b0;
assign COL[15156] = 1'b0;
assign COL[15157] = 1'b0;
assign COL[15158] = 1'b0;
assign COL[15159] = 1'b0;
assign COL[15160] = 1'b0;
assign COL[15161] = 1'b0;
assign COL[15162] = 1'b0;
assign COL[15163] = 1'b0;
assign COL[15164] = 1'b0;
assign COL[15165] = 1'b0;
assign COL[15166] = 1'b0;
assign COL[15167] = 1'b0;
assign COL[15168] = 1'b0;
assign COL[15169] = 1'b0;
assign COL[15170] = 1'b0;
assign COL[15171] = 1'b0;
assign COL[15172] = 1'b0;
assign COL[15173] = 1'b0;
assign COL[15174] = 1'b0;
assign COL[15175] = 1'b0;
assign COL[15176] = 1'b0;
assign COL[15177] = 1'b0;
assign COL[15178] = 1'b0;
assign COL[15179] = 1'b0;
assign COL[15180] = 1'b0;
assign COL[15181] = 1'b0;
assign COL[15182] = 1'b0;
assign COL[15183] = 1'b0;
assign COL[15184] = 1'b0;
assign COL[15185] = 1'b0;
assign COL[15186] = 1'b0;
assign COL[15187] = 1'b0;
assign COL[15188] = 1'b0;
assign COL[15189] = 1'b0;
assign COL[15190] = 1'b0;
assign COL[15191] = 1'b0;
assign COL[15192] = 1'b0;
assign COL[15193] = 1'b0;
assign COL[15194] = 1'b0;
assign COL[15195] = 1'b0;
assign COL[15196] = 1'b0;
assign COL[15197] = 1'b0;
assign COL[15198] = 1'b0;
assign COL[15199] = 1'b0;
assign COL[15200] = 1'b0;
assign COL[15201] = 1'b0;
assign COL[15202] = 1'b0;
assign COL[15203] = 1'b0;
assign COL[15204] = 1'b0;
assign COL[15205] = 1'b0;
assign COL[15206] = 1'b0;
assign COL[15207] = 1'b0;
assign COL[15208] = 1'b0;
assign COL[15209] = 1'b0;
assign COL[15210] = 1'b0;
assign COL[15211] = 1'b0;
assign COL[15212] = 1'b0;
assign COL[15213] = 1'b0;
assign COL[15214] = 1'b0;
assign COL[15215] = 1'b0;
assign COL[15216] = 1'b0;
assign COL[15217] = 1'b0;
assign COL[15218] = 1'b0;
assign COL[15219] = 1'b0;
assign COL[15220] = 1'b0;
assign COL[15221] = 1'b0;
assign COL[15222] = 1'b0;
assign COL[15223] = 1'b0;
assign COL[15224] = 1'b0;
assign COL[15225] = 1'b0;
assign COL[15226] = 1'b0;
assign COL[15227] = 1'b0;
assign COL[15228] = 1'b0;
assign COL[15229] = 1'b0;
assign COL[15230] = 1'b0;
assign COL[15231] = 1'b0;
assign COL[15232] = 1'b0;
assign COL[15233] = 1'b0;
assign COL[15234] = 1'b0;
assign COL[15235] = 1'b0;
assign COL[15236] = 1'b0;
assign COL[15237] = 1'b0;
assign COL[15238] = 1'b0;
assign COL[15239] = 1'b0;
assign COL[15240] = 1'b0;
assign COL[15241] = 1'b0;
assign COL[15242] = 1'b0;
assign COL[15243] = 1'b0;
assign COL[15244] = 1'b0;
assign COL[15245] = 1'b0;
assign COL[15246] = 1'b0;
assign COL[15247] = 1'b0;
assign COL[15248] = 1'b0;
assign COL[15249] = 1'b0;
assign COL[15250] = 1'b0;
assign COL[15251] = 1'b0;
assign COL[15252] = 1'b0;
assign COL[15253] = 1'b0;
assign COL[15254] = 1'b0;
assign COL[15255] = 1'b0;
assign COL[15256] = 1'b0;
assign COL[15257] = 1'b0;
assign COL[15258] = 1'b0;
assign COL[15259] = 1'b0;
assign COL[15260] = 1'b0;
assign COL[15261] = 1'b0;
assign COL[15262] = 1'b0;
assign COL[15263] = 1'b0;
assign COL[15264] = 1'b0;
assign COL[15265] = 1'b0;
assign COL[15266] = 1'b0;
assign COL[15267] = 1'b0;
assign COL[15268] = 1'b0;
assign COL[15269] = 1'b0;
assign COL[15270] = 1'b0;
assign COL[15271] = 1'b0;
assign COL[15272] = 1'b0;
assign COL[15273] = 1'b0;
assign COL[15274] = 1'b0;
assign COL[15275] = 1'b0;
assign COL[15276] = 1'b0;
assign COL[15277] = 1'b0;
assign COL[15278] = 1'b0;
assign COL[15279] = 1'b0;
assign COL[15280] = 1'b0;
assign COL[15281] = 1'b0;
assign COL[15282] = 1'b0;
assign COL[15283] = 1'b0;
assign COL[15284] = 1'b0;
assign COL[15285] = 1'b0;
assign COL[15286] = 1'b0;
assign COL[15287] = 1'b0;
assign COL[15288] = 1'b0;
assign COL[15289] = 1'b0;
assign COL[15290] = 1'b0;
assign COL[15291] = 1'b0;
assign COL[15292] = 1'b0;
assign COL[15293] = 1'b0;
assign COL[15294] = 1'b0;
assign COL[15295] = 1'b0;
assign COL[15296] = 1'b0;
assign COL[15297] = 1'b0;
assign COL[15298] = 1'b0;
assign COL[15299] = 1'b0;
assign COL[15300] = 1'b0;
assign COL[15301] = 1'b0;
assign COL[15302] = 1'b0;
assign COL[15303] = 1'b0;
assign COL[15304] = 1'b0;
assign COL[15305] = 1'b0;
assign COL[15306] = 1'b0;
assign COL[15307] = 1'b0;
assign COL[15308] = 1'b0;
assign COL[15309] = 1'b0;
assign COL[15310] = 1'b0;
assign COL[15311] = 1'b0;
assign COL[15312] = 1'b0;
assign COL[15313] = 1'b0;
assign COL[15314] = 1'b0;
assign COL[15315] = 1'b0;
assign COL[15316] = 1'b0;
assign COL[15317] = 1'b0;
assign COL[15318] = 1'b0;
assign COL[15319] = 1'b0;
assign COL[15320] = 1'b0;
assign COL[15321] = 1'b0;
assign COL[15322] = 1'b0;
assign COL[15323] = 1'b0;
assign COL[15324] = 1'b0;
assign COL[15325] = 1'b0;
assign COL[15326] = 1'b0;
assign COL[15327] = 1'b0;
assign COL[15328] = 1'b0;
assign COL[15329] = 1'b0;
assign COL[15330] = 1'b0;
assign COL[15331] = 1'b0;
assign COL[15332] = 1'b0;
assign COL[15333] = 1'b0;
assign COL[15334] = 1'b0;
assign COL[15335] = 1'b0;
assign COL[15336] = 1'b0;
assign COL[15337] = 1'b0;
assign COL[15338] = 1'b0;
assign COL[15339] = 1'b0;
assign COL[15340] = 1'b0;
assign COL[15341] = 1'b0;
assign COL[15342] = 1'b0;
assign COL[15343] = 1'b0;
assign COL[15344] = 1'b0;
assign COL[15345] = 1'b0;
assign COL[15346] = 1'b0;
assign COL[15347] = 1'b0;
assign COL[15348] = 1'b0;
assign COL[15349] = 1'b0;
assign COL[15350] = 1'b0;
assign COL[15351] = 1'b0;
assign COL[15352] = 1'b0;
assign COL[15353] = 1'b0;
assign COL[15354] = 1'b0;
assign COL[15355] = 1'b0;
assign COL[15356] = 1'b0;
assign COL[15357] = 1'b0;
assign COL[15358] = 1'b0;
assign COL[15359] = 1'b0;
assign COL[15360] = 1'b0;
assign COL[15361] = 1'b0;
assign COL[15362] = 1'b0;
assign COL[15363] = 1'b0;
assign COL[15364] = 1'b0;
assign COL[15365] = 1'b0;
assign COL[15366] = 1'b0;
assign COL[15367] = 1'b0;
assign COL[15368] = 1'b0;
assign COL[15369] = 1'b0;
assign COL[15370] = 1'b0;
assign COL[15371] = 1'b0;
assign COL[15372] = 1'b0;
assign COL[15373] = 1'b0;
assign COL[15374] = 1'b0;
assign COL[15375] = 1'b0;
assign COL[15376] = 1'b0;
assign COL[15377] = 1'b0;
assign COL[15378] = 1'b0;
assign COL[15379] = 1'b0;
assign COL[15380] = 1'b0;
assign COL[15381] = 1'b0;
assign COL[15382] = 1'b0;
assign COL[15383] = 1'b0;
assign COL[15384] = 1'b0;
assign COL[15385] = 1'b0;
assign COL[15386] = 1'b0;
assign COL[15387] = 1'b0;
assign COL[15388] = 1'b0;
assign COL[15389] = 1'b0;
assign COL[15390] = 1'b0;
assign COL[15391] = 1'b0;
assign COL[15392] = 1'b0;
assign COL[15393] = 1'b0;
assign COL[15394] = 1'b0;
assign COL[15395] = 1'b0;
assign COL[15396] = 1'b0;
assign COL[15397] = 1'b0;
assign COL[15398] = 1'b0;
assign COL[15399] = 1'b0;
assign COL[15400] = 1'b0;
assign COL[15401] = 1'b0;
assign COL[15402] = 1'b0;
assign COL[15403] = 1'b0;
assign COL[15404] = 1'b0;
assign COL[15405] = 1'b0;
assign COL[15406] = 1'b0;
assign COL[15407] = 1'b0;
assign COL[15408] = 1'b0;
assign COL[15409] = 1'b0;
assign COL[15410] = 1'b0;
assign COL[15411] = 1'b0;
assign COL[15412] = 1'b0;
assign COL[15413] = 1'b0;
assign COL[15414] = 1'b0;
assign COL[15415] = 1'b0;
assign COL[15416] = 1'b0;
assign COL[15417] = 1'b0;
assign COL[15418] = 1'b0;
assign COL[15419] = 1'b0;
assign COL[15420] = 1'b0;
assign COL[15421] = 1'b0;
assign COL[15422] = 1'b0;
assign COL[15423] = 1'b0;
assign COL[15424] = 1'b0;
assign COL[15425] = 1'b0;
assign COL[15426] = 1'b0;
assign COL[15427] = 1'b0;
assign COL[15428] = 1'b0;
assign COL[15429] = 1'b0;
assign COL[15430] = 1'b0;
assign COL[15431] = 1'b0;
assign COL[15432] = 1'b0;
assign COL[15433] = 1'b0;
assign COL[15434] = 1'b0;
assign COL[15435] = 1'b0;
assign COL[15436] = 1'b0;
assign COL[15437] = 1'b0;
assign COL[15438] = 1'b0;
assign COL[15439] = 1'b0;
assign COL[15440] = 1'b0;
assign COL[15441] = 1'b0;
assign COL[15442] = 1'b0;
assign COL[15443] = 1'b0;
assign COL[15444] = 1'b0;
assign COL[15445] = 1'b0;
assign COL[15446] = 1'b0;
assign COL[15447] = 1'b0;
assign COL[15448] = 1'b0;
assign COL[15449] = 1'b0;
assign COL[15450] = 1'b0;
assign COL[15451] = 1'b0;
assign COL[15452] = 1'b0;
assign COL[15453] = 1'b0;
assign COL[15454] = 1'b0;
assign COL[15455] = 1'b0;
assign COL[15456] = 1'b0;
assign COL[15457] = 1'b0;
assign COL[15458] = 1'b0;
assign COL[15459] = 1'b0;
assign COL[15460] = 1'b0;
assign COL[15461] = 1'b0;
assign COL[15462] = 1'b0;
assign COL[15463] = 1'b0;
assign COL[15464] = 1'b0;
assign COL[15465] = 1'b0;
assign COL[15466] = 1'b0;
assign COL[15467] = 1'b0;
assign COL[15468] = 1'b0;
assign COL[15469] = 1'b0;
assign COL[15470] = 1'b0;
assign COL[15471] = 1'b0;
assign COL[15472] = 1'b0;
assign COL[15473] = 1'b0;
assign COL[15474] = 1'b0;
assign COL[15475] = 1'b0;
assign COL[15476] = 1'b0;
assign COL[15477] = 1'b0;
assign COL[15478] = 1'b0;
assign COL[15479] = 1'b0;
assign COL[15480] = 1'b0;
assign COL[15481] = 1'b0;
assign COL[15482] = 1'b0;
assign COL[15483] = 1'b0;
assign COL[15484] = 1'b0;
assign COL[15485] = 1'b0;
assign COL[15486] = 1'b0;
assign COL[15487] = 1'b0;
assign COL[15488] = 1'b0;
assign COL[15489] = 1'b0;
assign COL[15490] = 1'b0;
assign COL[15491] = 1'b0;
assign COL[15492] = 1'b0;
assign COL[15493] = 1'b0;
assign COL[15494] = 1'b0;
assign COL[15495] = 1'b0;
assign COL[15496] = 1'b0;
assign COL[15497] = 1'b0;
assign COL[15498] = 1'b0;
assign COL[15499] = 1'b0;
assign COL[15500] = 1'b0;
assign COL[15501] = 1'b0;
assign COL[15502] = 1'b0;
assign COL[15503] = 1'b0;
assign COL[15504] = 1'b0;
assign COL[15505] = 1'b0;
assign COL[15506] = 1'b0;
assign COL[15507] = 1'b0;
assign COL[15508] = 1'b0;
assign COL[15509] = 1'b0;
assign COL[15510] = 1'b0;
assign COL[15511] = 1'b0;
assign COL[15512] = 1'b0;
assign COL[15513] = 1'b0;
assign COL[15514] = 1'b0;
assign COL[15515] = 1'b0;
assign COL[15516] = 1'b0;
assign COL[15517] = 1'b0;
assign COL[15518] = 1'b0;
assign COL[15519] = 1'b0;
assign COL[15520] = 1'b0;
assign COL[15521] = 1'b0;
assign COL[15522] = 1'b0;
assign COL[15523] = 1'b0;
assign COL[15524] = 1'b0;
assign COL[15525] = 1'b0;
assign COL[15526] = 1'b0;
assign COL[15527] = 1'b0;
assign COL[15528] = 1'b0;
assign COL[15529] = 1'b0;
assign COL[15530] = 1'b0;
assign COL[15531] = 1'b0;
assign COL[15532] = 1'b0;
assign COL[15533] = 1'b0;
assign COL[15534] = 1'b0;
assign COL[15535] = 1'b0;
assign COL[15536] = 1'b0;
assign COL[15537] = 1'b0;
assign COL[15538] = 1'b0;
assign COL[15539] = 1'b0;
assign COL[15540] = 1'b0;
assign COL[15541] = 1'b0;
assign COL[15542] = 1'b0;
assign COL[15543] = 1'b0;
assign COL[15544] = 1'b0;
assign COL[15545] = 1'b0;
assign COL[15546] = 1'b0;
assign COL[15547] = 1'b0;
assign COL[15548] = 1'b0;
assign COL[15549] = 1'b0;
assign COL[15550] = 1'b0;
assign COL[15551] = 1'b0;
assign COL[15552] = 1'b0;
assign COL[15553] = 1'b0;
assign COL[15554] = 1'b0;
assign COL[15555] = 1'b0;
assign COL[15556] = 1'b0;
assign COL[15557] = 1'b0;
assign COL[15558] = 1'b0;
assign COL[15559] = 1'b0;
assign COL[15560] = 1'b0;
assign COL[15561] = 1'b0;
assign COL[15562] = 1'b0;
assign COL[15563] = 1'b0;
assign COL[15564] = 1'b0;
assign COL[15565] = 1'b0;
assign COL[15566] = 1'b0;
assign COL[15567] = 1'b0;
assign COL[15568] = 1'b0;
assign COL[15569] = 1'b0;
assign COL[15570] = 1'b0;
assign COL[15571] = 1'b0;
assign COL[15572] = 1'b0;
assign COL[15573] = 1'b0;
assign COL[15574] = 1'b0;
assign COL[15575] = 1'b0;
assign COL[15576] = 1'b0;
assign COL[15577] = 1'b0;
assign COL[15578] = 1'b0;
assign COL[15579] = 1'b0;
assign COL[15580] = 1'b0;
assign COL[15581] = 1'b0;
assign COL[15582] = 1'b0;
assign COL[15583] = 1'b0;
assign COL[15584] = 1'b0;
assign COL[15585] = 1'b0;
assign COL[15586] = 1'b0;
assign COL[15587] = 1'b0;
assign COL[15588] = 1'b0;
assign COL[15589] = 1'b0;
assign COL[15590] = 1'b0;
assign COL[15591] = 1'b0;
assign COL[15592] = 1'b0;
assign COL[15593] = 1'b0;
assign COL[15594] = 1'b0;
assign COL[15595] = 1'b0;
assign COL[15596] = 1'b0;
assign COL[15597] = 1'b0;
assign COL[15598] = 1'b0;
assign COL[15599] = 1'b0;
assign COL[15600] = 1'b0;
assign COL[15601] = 1'b0;
assign COL[15602] = 1'b0;
assign COL[15603] = 1'b0;
assign COL[15604] = 1'b0;
assign COL[15605] = 1'b0;
assign COL[15606] = 1'b0;
assign COL[15607] = 1'b0;
assign COL[15608] = 1'b0;
assign COL[15609] = 1'b0;
assign COL[15610] = 1'b0;
assign COL[15611] = 1'b0;
assign COL[15612] = 1'b0;
assign COL[15613] = 1'b0;
assign COL[15614] = 1'b0;
assign COL[15615] = 1'b0;
assign COL[15616] = 1'b0;
assign COL[15617] = 1'b0;
assign COL[15618] = 1'b0;
assign COL[15619] = 1'b0;
assign COL[15620] = 1'b0;
assign COL[15621] = 1'b0;
assign COL[15622] = 1'b0;
assign COL[15623] = 1'b0;
assign COL[15624] = 1'b0;
assign COL[15625] = 1'b0;
assign COL[15626] = 1'b0;
assign COL[15627] = 1'b0;
assign COL[15628] = 1'b0;
assign COL[15629] = 1'b0;
assign COL[15630] = 1'b0;
assign COL[15631] = 1'b0;
assign COL[15632] = 1'b0;
assign COL[15633] = 1'b0;
assign COL[15634] = 1'b0;
assign COL[15635] = 1'b0;
assign COL[15636] = 1'b0;
assign COL[15637] = 1'b0;
assign COL[15638] = 1'b0;
assign COL[15639] = 1'b0;
assign COL[15640] = 1'b0;
assign COL[15641] = 1'b0;
assign COL[15642] = 1'b0;
assign COL[15643] = 1'b0;
assign COL[15644] = 1'b0;
assign COL[15645] = 1'b0;
assign COL[15646] = 1'b0;
assign COL[15647] = 1'b0;
assign COL[15648] = 1'b0;
assign COL[15649] = 1'b0;
assign COL[15650] = 1'b0;
assign COL[15651] = 1'b0;
assign COL[15652] = 1'b0;
assign COL[15653] = 1'b0;
assign COL[15654] = 1'b0;
assign COL[15655] = 1'b0;
assign COL[15656] = 1'b0;
assign COL[15657] = 1'b0;
assign COL[15658] = 1'b0;
assign COL[15659] = 1'b0;
assign COL[15660] = 1'b0;
assign COL[15661] = 1'b0;
assign COL[15662] = 1'b0;
assign COL[15663] = 1'b0;
assign COL[15664] = 1'b0;
assign COL[15665] = 1'b0;
assign COL[15666] = 1'b0;
assign COL[15667] = 1'b0;
assign COL[15668] = 1'b0;
assign COL[15669] = 1'b0;
assign COL[15670] = 1'b0;
assign COL[15671] = 1'b0;
assign COL[15672] = 1'b0;
assign COL[15673] = 1'b0;
assign COL[15674] = 1'b0;
assign COL[15675] = 1'b0;
assign COL[15676] = 1'b0;
assign COL[15677] = 1'b0;
assign COL[15678] = 1'b0;
assign COL[15679] = 1'b0;
assign COL[15680] = 1'b0;
assign COL[15681] = 1'b0;
assign COL[15682] = 1'b0;
assign COL[15683] = 1'b0;
assign COL[15684] = 1'b0;
assign COL[15685] = 1'b0;
assign COL[15686] = 1'b0;
assign COL[15687] = 1'b0;
assign COL[15688] = 1'b0;
assign COL[15689] = 1'b0;
assign COL[15690] = 1'b0;
assign COL[15691] = 1'b0;
assign COL[15692] = 1'b0;
assign COL[15693] = 1'b0;
assign COL[15694] = 1'b0;
assign COL[15695] = 1'b0;
assign COL[15696] = 1'b0;
assign COL[15697] = 1'b0;
assign COL[15698] = 1'b0;
assign COL[15699] = 1'b0;
assign COL[15700] = 1'b0;
assign COL[15701] = 1'b0;
assign COL[15702] = 1'b0;
assign COL[15703] = 1'b0;
assign COL[15704] = 1'b0;
assign COL[15705] = 1'b0;
assign COL[15706] = 1'b0;
assign COL[15707] = 1'b0;
assign COL[15708] = 1'b0;
assign COL[15709] = 1'b0;
assign COL[15710] = 1'b0;
assign COL[15711] = 1'b0;
assign COL[15712] = 1'b0;
assign COL[15713] = 1'b0;
assign COL[15714] = 1'b0;
assign COL[15715] = 1'b0;
assign COL[15716] = 1'b0;
assign COL[15717] = 1'b0;
assign COL[15718] = 1'b0;
assign COL[15719] = 1'b0;
assign COL[15720] = 1'b0;
assign COL[15721] = 1'b0;
assign COL[15722] = 1'b0;
assign COL[15723] = 1'b0;
assign COL[15724] = 1'b0;
assign COL[15725] = 1'b0;
assign COL[15726] = 1'b0;
assign COL[15727] = 1'b0;
assign COL[15728] = 1'b0;
assign COL[15729] = 1'b0;
assign COL[15730] = 1'b0;
assign COL[15731] = 1'b0;
assign COL[15732] = 1'b0;
assign COL[15733] = 1'b0;
assign COL[15734] = 1'b0;
assign COL[15735] = 1'b0;
assign COL[15736] = 1'b0;
assign COL[15737] = 1'b0;
assign COL[15738] = 1'b0;
assign COL[15739] = 1'b0;
assign COL[15740] = 1'b0;
assign COL[15741] = 1'b0;
assign COL[15742] = 1'b0;
assign COL[15743] = 1'b0;
assign COL[15744] = 1'b0;
assign COL[15745] = 1'b0;
assign COL[15746] = 1'b0;
assign COL[15747] = 1'b0;
assign COL[15748] = 1'b0;
assign COL[15749] = 1'b0;
assign COL[15750] = 1'b0;
assign COL[15751] = 1'b0;
assign COL[15752] = 1'b0;
assign COL[15753] = 1'b0;
assign COL[15754] = 1'b0;
assign COL[15755] = 1'b0;
assign COL[15756] = 1'b0;
assign COL[15757] = 1'b0;
assign COL[15758] = 1'b0;
assign COL[15759] = 1'b0;
assign COL[15760] = 1'b0;
assign COL[15761] = 1'b0;
assign COL[15762] = 1'b0;
assign COL[15763] = 1'b0;
assign COL[15764] = 1'b0;
assign COL[15765] = 1'b0;
assign COL[15766] = 1'b0;
assign COL[15767] = 1'b0;
assign COL[15768] = 1'b0;
assign COL[15769] = 1'b0;
assign COL[15770] = 1'b0;
assign COL[15771] = 1'b0;
assign COL[15772] = 1'b0;
assign COL[15773] = 1'b0;
assign COL[15774] = 1'b0;
assign COL[15775] = 1'b0;
assign COL[15776] = 1'b0;
assign COL[15777] = 1'b0;
assign COL[15778] = 1'b0;
assign COL[15779] = 1'b0;
assign COL[15780] = 1'b0;
assign COL[15781] = 1'b0;
assign COL[15782] = 1'b0;
assign COL[15783] = 1'b0;
assign COL[15784] = 1'b0;
assign COL[15785] = 1'b0;
assign COL[15786] = 1'b0;
assign COL[15787] = 1'b0;
assign COL[15788] = 1'b0;
assign COL[15789] = 1'b0;
assign COL[15790] = 1'b0;
assign COL[15791] = 1'b0;
assign COL[15792] = 1'b0;
assign COL[15793] = 1'b0;
assign COL[15794] = 1'b0;
assign COL[15795] = 1'b0;
assign COL[15796] = 1'b0;
assign COL[15797] = 1'b0;
assign COL[15798] = 1'b0;
assign COL[15799] = 1'b0;
assign COL[15800] = 1'b0;
assign COL[15801] = 1'b0;
assign COL[15802] = 1'b0;
assign COL[15803] = 1'b0;
assign COL[15804] = 1'b0;
assign COL[15805] = 1'b0;
assign COL[15806] = 1'b0;
assign COL[15807] = 1'b0;
assign COL[15808] = 1'b0;
assign COL[15809] = 1'b0;
assign COL[15810] = 1'b0;
assign COL[15811] = 1'b0;
assign COL[15812] = 1'b0;
assign COL[15813] = 1'b0;
assign COL[15814] = 1'b0;
assign COL[15815] = 1'b0;
assign COL[15816] = 1'b0;
assign COL[15817] = 1'b0;
assign COL[15818] = 1'b0;
assign COL[15819] = 1'b0;
assign COL[15820] = 1'b0;
assign COL[15821] = 1'b0;
assign COL[15822] = 1'b0;
assign COL[15823] = 1'b0;
assign COL[15824] = 1'b0;
assign COL[15825] = 1'b0;
assign COL[15826] = 1'b0;
assign COL[15827] = 1'b0;
assign COL[15828] = 1'b0;
assign COL[15829] = 1'b0;
assign COL[15830] = 1'b0;
assign COL[15831] = 1'b0;
assign COL[15832] = 1'b0;
assign COL[15833] = 1'b0;
assign COL[15834] = 1'b0;
assign COL[15835] = 1'b0;
assign COL[15836] = 1'b0;
assign COL[15837] = 1'b0;
assign COL[15838] = 1'b0;
assign COL[15839] = 1'b0;
assign COL[15840] = 1'b0;
assign COL[15841] = 1'b0;
assign COL[15842] = 1'b0;
assign COL[15843] = 1'b0;
assign COL[15844] = 1'b0;
assign COL[15845] = 1'b0;
assign COL[15846] = 1'b0;
assign COL[15847] = 1'b0;
assign COL[15848] = 1'b0;
assign COL[15849] = 1'b0;
assign COL[15850] = 1'b0;
assign COL[15851] = 1'b0;
assign COL[15852] = 1'b0;
assign COL[15853] = 1'b0;
assign COL[15854] = 1'b0;
assign COL[15855] = 1'b0;
assign COL[15856] = 1'b0;
assign COL[15857] = 1'b0;
assign COL[15858] = 1'b0;
assign COL[15859] = 1'b0;
assign COL[15860] = 1'b0;
assign COL[15861] = 1'b0;
assign COL[15862] = 1'b0;
assign COL[15863] = 1'b0;
assign COL[15864] = 1'b0;
assign COL[15865] = 1'b0;
assign COL[15866] = 1'b0;
assign COL[15867] = 1'b0;
assign COL[15868] = 1'b0;
assign COL[15869] = 1'b0;
assign COL[15870] = 1'b0;
assign COL[15871] = 1'b0;
assign COL[15872] = 1'b0;
assign COL[15873] = 1'b0;
assign COL[15874] = 1'b0;
assign COL[15875] = 1'b0;
assign COL[15876] = 1'b0;
assign COL[15877] = 1'b0;
assign COL[15878] = 1'b0;
assign COL[15879] = 1'b0;
assign COL[15880] = 1'b0;
assign COL[15881] = 1'b0;
assign COL[15882] = 1'b0;
assign COL[15883] = 1'b0;
assign COL[15884] = 1'b0;
assign COL[15885] = 1'b0;
assign COL[15886] = 1'b0;
assign COL[15887] = 1'b0;
assign COL[15888] = 1'b0;
assign COL[15889] = 1'b0;
assign COL[15890] = 1'b0;
assign COL[15891] = 1'b0;
assign COL[15892] = 1'b0;
assign COL[15893] = 1'b0;
assign COL[15894] = 1'b0;
assign COL[15895] = 1'b0;
assign COL[15896] = 1'b0;
assign COL[15897] = 1'b0;
assign COL[15898] = 1'b0;
assign COL[15899] = 1'b0;
assign COL[15900] = 1'b0;
assign COL[15901] = 1'b0;
assign COL[15902] = 1'b0;
assign COL[15903] = 1'b0;
assign COL[15904] = 1'b0;
assign COL[15905] = 1'b0;
assign COL[15906] = 1'b0;
assign COL[15907] = 1'b0;
assign COL[15908] = 1'b0;
assign COL[15909] = 1'b0;
assign COL[15910] = 1'b0;
assign COL[15911] = 1'b0;
assign COL[15912] = 1'b0;
assign COL[15913] = 1'b0;
assign COL[15914] = 1'b0;
assign COL[15915] = 1'b0;
assign COL[15916] = 1'b0;
assign COL[15917] = 1'b0;
assign COL[15918] = 1'b0;
assign COL[15919] = 1'b0;
assign COL[15920] = 1'b0;
assign COL[15921] = 1'b0;
assign COL[15922] = 1'b0;
assign COL[15923] = 1'b0;
assign COL[15924] = 1'b0;
assign COL[15925] = 1'b0;
assign COL[15926] = 1'b0;
assign COL[15927] = 1'b0;
assign COL[15928] = 1'b0;
assign COL[15929] = 1'b0;
assign COL[15930] = 1'b0;
assign COL[15931] = 1'b0;
assign COL[15932] = 1'b0;
assign COL[15933] = 1'b0;
assign COL[15934] = 1'b0;
assign COL[15935] = 1'b0;
assign COL[15936] = 1'b0;
assign COL[15937] = 1'b0;
assign COL[15938] = 1'b0;
assign COL[15939] = 1'b0;
assign COL[15940] = 1'b0;
assign COL[15941] = 1'b0;
assign COL[15942] = 1'b0;
assign COL[15943] = 1'b0;
assign COL[15944] = 1'b0;
assign COL[15945] = 1'b0;
assign COL[15946] = 1'b0;
assign COL[15947] = 1'b0;
assign COL[15948] = 1'b0;
assign COL[15949] = 1'b0;
assign COL[15950] = 1'b0;
assign COL[15951] = 1'b0;
assign COL[15952] = 1'b0;
assign COL[15953] = 1'b0;
assign COL[15954] = 1'b0;
assign COL[15955] = 1'b0;
assign COL[15956] = 1'b0;
assign COL[15957] = 1'b0;
assign COL[15958] = 1'b0;
assign COL[15959] = 1'b0;
assign COL[15960] = 1'b0;
assign COL[15961] = 1'b0;
assign COL[15962] = 1'b0;
assign COL[15963] = 1'b0;
assign COL[15964] = 1'b0;
assign COL[15965] = 1'b0;
assign COL[15966] = 1'b0;
assign COL[15967] = 1'b0;
assign COL[15968] = 1'b0;
assign COL[15969] = 1'b0;
assign COL[15970] = 1'b0;
assign COL[15971] = 1'b0;
assign COL[15972] = 1'b0;
assign COL[15973] = 1'b0;
assign COL[15974] = 1'b0;
assign COL[15975] = 1'b0;
assign COL[15976] = 1'b0;
assign COL[15977] = 1'b0;
assign COL[15978] = 1'b0;
assign COL[15979] = 1'b0;
assign COL[15980] = 1'b0;
assign COL[15981] = 1'b0;
assign COL[15982] = 1'b0;
assign COL[15983] = 1'b0;
assign COL[15984] = 1'b0;
assign COL[15985] = 1'b0;
assign COL[15986] = 1'b0;
assign COL[15987] = 1'b0;
assign COL[15988] = 1'b0;
assign COL[15989] = 1'b0;
assign COL[15990] = 1'b0;
assign COL[15991] = 1'b0;
assign COL[15992] = 1'b0;
assign COL[15993] = 1'b0;
assign COL[15994] = 1'b0;
assign COL[15995] = 1'b0;
assign COL[15996] = 1'b0;
assign COL[15997] = 1'b0;
assign COL[15998] = 1'b0;
assign COL[15999] = 1'b0;
assign COL[16000] = 1'b0;
assign COL[16001] = 1'b0;
assign COL[16002] = 1'b0;
assign COL[16003] = 1'b0;
assign COL[16004] = 1'b0;
assign COL[16005] = 1'b0;
assign COL[16006] = 1'b0;
assign COL[16007] = 1'b0;
assign COL[16008] = 1'b0;
assign COL[16009] = 1'b0;
assign COL[16010] = 1'b0;
assign COL[16011] = 1'b0;
assign COL[16012] = 1'b0;
assign COL[16013] = 1'b0;
assign COL[16014] = 1'b0;
assign COL[16015] = 1'b0;
assign COL[16016] = 1'b0;
assign COL[16017] = 1'b0;
assign COL[16018] = 1'b0;
assign COL[16019] = 1'b0;
assign COL[16020] = 1'b0;
assign COL[16021] = 1'b0;
assign COL[16022] = 1'b0;
assign COL[16023] = 1'b0;
assign COL[16024] = 1'b0;
assign COL[16025] = 1'b0;
assign COL[16026] = 1'b0;
assign COL[16027] = 1'b0;
assign COL[16028] = 1'b0;
assign COL[16029] = 1'b0;
assign COL[16030] = 1'b0;
assign COL[16031] = 1'b0;
assign COL[16032] = 1'b0;
assign COL[16033] = 1'b0;
assign COL[16034] = 1'b0;
assign COL[16035] = 1'b0;
assign COL[16036] = 1'b0;
assign COL[16037] = 1'b0;
assign COL[16038] = 1'b0;
assign COL[16039] = 1'b0;
assign COL[16040] = 1'b0;
assign COL[16041] = 1'b0;
assign COL[16042] = 1'b0;
assign COL[16043] = 1'b0;
assign COL[16044] = 1'b0;
assign COL[16045] = 1'b0;
assign COL[16046] = 1'b0;
assign COL[16047] = 1'b0;
assign COL[16048] = 1'b0;
assign COL[16049] = 1'b0;
assign COL[16050] = 1'b0;
assign COL[16051] = 1'b0;
assign COL[16052] = 1'b0;
assign COL[16053] = 1'b0;
assign COL[16054] = 1'b0;
assign COL[16055] = 1'b0;
assign COL[16056] = 1'b0;
assign COL[16057] = 1'b0;
assign COL[16058] = 1'b0;
assign COL[16059] = 1'b0;
assign COL[16060] = 1'b0;
assign COL[16061] = 1'b0;
assign COL[16062] = 1'b0;
assign COL[16063] = 1'b0;
assign COL[16064] = 1'b0;
assign COL[16065] = 1'b0;
assign COL[16066] = 1'b0;
assign COL[16067] = 1'b0;
assign COL[16068] = 1'b0;
assign COL[16069] = 1'b0;
assign COL[16070] = 1'b0;
assign COL[16071] = 1'b0;
assign COL[16072] = 1'b0;
assign COL[16073] = 1'b0;
assign COL[16074] = 1'b0;
assign COL[16075] = 1'b0;
assign COL[16076] = 1'b0;
assign COL[16077] = 1'b0;
assign COL[16078] = 1'b0;
assign COL[16079] = 1'b0;
assign COL[16080] = 1'b0;
assign COL[16081] = 1'b0;
assign COL[16082] = 1'b0;
assign COL[16083] = 1'b0;
assign COL[16084] = 1'b0;
assign COL[16085] = 1'b0;
assign COL[16086] = 1'b0;
assign COL[16087] = 1'b0;
assign COL[16088] = 1'b0;
assign COL[16089] = 1'b0;
assign COL[16090] = 1'b0;
assign COL[16091] = 1'b0;
assign COL[16092] = 1'b0;
assign COL[16093] = 1'b0;
assign COL[16094] = 1'b0;
assign COL[16095] = 1'b0;
assign COL[16096] = 1'b0;
assign COL[16097] = 1'b0;
assign COL[16098] = 1'b0;
assign COL[16099] = 1'b0;
assign COL[16100] = 1'b0;
assign COL[16101] = 1'b0;
assign COL[16102] = 1'b0;
assign COL[16103] = 1'b0;
assign COL[16104] = 1'b0;
assign COL[16105] = 1'b0;
assign COL[16106] = 1'b0;
assign COL[16107] = 1'b0;
assign COL[16108] = 1'b0;
assign COL[16109] = 1'b0;
assign COL[16110] = 1'b0;
assign COL[16111] = 1'b0;
assign COL[16112] = 1'b0;
assign COL[16113] = 1'b0;
assign COL[16114] = 1'b0;
assign COL[16115] = 1'b0;
assign COL[16116] = 1'b0;
assign COL[16117] = 1'b0;
assign COL[16118] = 1'b0;
assign COL[16119] = 1'b0;
assign COL[16120] = 1'b0;
assign COL[16121] = 1'b0;
assign COL[16122] = 1'b0;
assign COL[16123] = 1'b0;
assign COL[16124] = 1'b0;
assign COL[16125] = 1'b0;
assign COL[16126] = 1'b0;
assign COL[16127] = 1'b0;
assign COL[16128] = 1'b0;
assign COL[16129] = 1'b0;
assign COL[16130] = 1'b0;
assign COL[16131] = 1'b0;
assign COL[16132] = 1'b0;
assign COL[16133] = 1'b0;
assign COL[16134] = 1'b0;
assign COL[16135] = 1'b0;
assign COL[16136] = 1'b0;
assign COL[16137] = 1'b0;
assign COL[16138] = 1'b0;
assign COL[16139] = 1'b0;
assign COL[16140] = 1'b0;
assign COL[16141] = 1'b0;
assign COL[16142] = 1'b0;
assign COL[16143] = 1'b0;
assign COL[16144] = 1'b0;
assign COL[16145] = 1'b0;
assign COL[16146] = 1'b0;
assign COL[16147] = 1'b0;
assign COL[16148] = 1'b0;
assign COL[16149] = 1'b0;
assign COL[16150] = 1'b0;
assign COL[16151] = 1'b0;
assign COL[16152] = 1'b0;
assign COL[16153] = 1'b0;
assign COL[16154] = 1'b0;
assign COL[16155] = 1'b0;
assign COL[16156] = 1'b0;
assign COL[16157] = 1'b0;
assign COL[16158] = 1'b0;
assign COL[16159] = 1'b0;
assign COL[16160] = 1'b0;
assign COL[16161] = 1'b0;
assign COL[16162] = 1'b0;
assign COL[16163] = 1'b0;
assign COL[16164] = 1'b0;
assign COL[16165] = 1'b0;
assign COL[16166] = 1'b0;
assign COL[16167] = 1'b0;
assign COL[16168] = 1'b0;
assign COL[16169] = 1'b0;
assign COL[16170] = 1'b0;
assign COL[16171] = 1'b0;
assign COL[16172] = 1'b0;
assign COL[16173] = 1'b0;
assign COL[16174] = 1'b0;
assign COL[16175] = 1'b0;
assign COL[16176] = 1'b0;
assign COL[16177] = 1'b0;
assign COL[16178] = 1'b0;
assign COL[16179] = 1'b0;
assign COL[16180] = 1'b0;
assign COL[16181] = 1'b0;
assign COL[16182] = 1'b0;
assign COL[16183] = 1'b0;
assign COL[16184] = 1'b0;
assign COL[16185] = 1'b0;
assign COL[16186] = 1'b0;
assign COL[16187] = 1'b0;
assign COL[16188] = 1'b0;
assign COL[16189] = 1'b0;
assign COL[16190] = 1'b0;
assign COL[16191] = 1'b0;
assign COL[16192] = 1'b0;
assign COL[16193] = 1'b0;
assign COL[16194] = 1'b0;
assign COL[16195] = 1'b0;
assign COL[16196] = 1'b0;
assign COL[16197] = 1'b0;
assign COL[16198] = 1'b0;
assign COL[16199] = 1'b0;
assign COL[16200] = 1'b0;
assign COL[16201] = 1'b0;
assign COL[16202] = 1'b0;
assign COL[16203] = 1'b0;
assign COL[16204] = 1'b0;
assign COL[16205] = 1'b0;
assign COL[16206] = 1'b0;
assign COL[16207] = 1'b0;
assign COL[16208] = 1'b0;
assign COL[16209] = 1'b0;
assign COL[16210] = 1'b0;
assign COL[16211] = 1'b0;
assign COL[16212] = 1'b0;
assign COL[16213] = 1'b0;
assign COL[16214] = 1'b0;
assign COL[16215] = 1'b0;
assign COL[16216] = 1'b0;
assign COL[16217] = 1'b0;
assign COL[16218] = 1'b0;
assign COL[16219] = 1'b0;
assign COL[16220] = 1'b0;
assign COL[16221] = 1'b0;
assign COL[16222] = 1'b0;
assign COL[16223] = 1'b0;
assign COL[16224] = 1'b0;
assign COL[16225] = 1'b0;
assign COL[16226] = 1'b0;
assign COL[16227] = 1'b0;
assign COL[16228] = 1'b0;
assign COL[16229] = 1'b0;
assign COL[16230] = 1'b0;
assign COL[16231] = 1'b0;
assign COL[16232] = 1'b0;
assign COL[16233] = 1'b0;
assign COL[16234] = 1'b0;
assign COL[16235] = 1'b0;
assign COL[16236] = 1'b0;
assign COL[16237] = 1'b0;
assign COL[16238] = 1'b0;
assign COL[16239] = 1'b0;
assign COL[16240] = 1'b0;
assign COL[16241] = 1'b0;
assign COL[16242] = 1'b0;
assign COL[16243] = 1'b0;
assign COL[16244] = 1'b0;
assign COL[16245] = 1'b0;
assign COL[16246] = 1'b0;
assign COL[16247] = 1'b0;
assign COL[16248] = 1'b0;
assign COL[16249] = 1'b0;
assign COL[16250] = 1'b0;
assign COL[16251] = 1'b0;
assign COL[16252] = 1'b0;
assign COL[16253] = 1'b0;
assign COL[16254] = 1'b0;
assign COL[16255] = 1'b0;
assign COL[16256] = 1'b0;
assign COL[16257] = 1'b0;
assign COL[16258] = 1'b0;
assign COL[16259] = 1'b0;
assign COL[16260] = 1'b0;
assign COL[16261] = 1'b0;
assign COL[16262] = 1'b0;
assign COL[16263] = 1'b0;
assign COL[16264] = 1'b0;
assign COL[16265] = 1'b0;
assign COL[16266] = 1'b0;
assign COL[16267] = 1'b0;
assign COL[16268] = 1'b0;
assign COL[16269] = 1'b0;
assign COL[16270] = 1'b0;
assign COL[16271] = 1'b0;
assign COL[16272] = 1'b0;
assign COL[16273] = 1'b0;
assign COL[16274] = 1'b0;
assign COL[16275] = 1'b0;
assign COL[16276] = 1'b0;
assign COL[16277] = 1'b0;
assign COL[16278] = 1'b0;
assign COL[16279] = 1'b0;
assign COL[16280] = 1'b0;
assign COL[16281] = 1'b0;
assign COL[16282] = 1'b0;
assign COL[16283] = 1'b0;
assign COL[16284] = 1'b0;
assign COL[16285] = 1'b0;
assign COL[16286] = 1'b0;
assign COL[16287] = 1'b0;
assign COL[16288] = 1'b0;
assign COL[16289] = 1'b0;
assign COL[16290] = 1'b0;
assign COL[16291] = 1'b0;
assign COL[16292] = 1'b0;
assign COL[16293] = 1'b0;
assign COL[16294] = 1'b0;
assign COL[16295] = 1'b0;
assign COL[16296] = 1'b0;
assign COL[16297] = 1'b0;
assign COL[16298] = 1'b0;
assign COL[16299] = 1'b0;
assign COL[16300] = 1'b0;
assign COL[16301] = 1'b0;
assign COL[16302] = 1'b0;
assign COL[16303] = 1'b0;
assign COL[16304] = 1'b0;
assign COL[16305] = 1'b0;
assign COL[16306] = 1'b0;
assign COL[16307] = 1'b0;
assign COL[16308] = 1'b0;
assign COL[16309] = 1'b0;
assign COL[16310] = 1'b0;
assign COL[16311] = 1'b0;
assign COL[16312] = 1'b0;
assign COL[16313] = 1'b0;
assign COL[16314] = 1'b0;
assign COL[16315] = 1'b0;
assign COL[16316] = 1'b0;
assign COL[16317] = 1'b0;
assign COL[16318] = 1'b0;
assign COL[16319] = 1'b0;
assign COL[16320] = 1'b0;
assign COL[16321] = 1'b0;
assign COL[16322] = 1'b0;
assign COL[16323] = 1'b0;
assign COL[16324] = 1'b0;
assign COL[16325] = 1'b0;
assign COL[16326] = 1'b0;
assign COL[16327] = 1'b0;
assign COL[16328] = 1'b0;
assign COL[16329] = 1'b0;
assign COL[16330] = 1'b0;
assign COL[16331] = 1'b0;
assign COL[16332] = 1'b0;
assign COL[16333] = 1'b0;
assign COL[16334] = 1'b0;
assign COL[16335] = 1'b0;
assign COL[16336] = 1'b0;
assign COL[16337] = 1'b0;
assign COL[16338] = 1'b0;
assign COL[16339] = 1'b0;
assign COL[16340] = 1'b0;
assign COL[16341] = 1'b0;
assign COL[16342] = 1'b0;
assign COL[16343] = 1'b0;
assign COL[16344] = 1'b0;
assign COL[16345] = 1'b0;
assign COL[16346] = 1'b0;
assign COL[16347] = 1'b0;
assign COL[16348] = 1'b0;
assign COL[16349] = 1'b0;
assign COL[16350] = 1'b0;
assign COL[16351] = 1'b0;
assign COL[16352] = 1'b0;
assign COL[16353] = 1'b0;
assign COL[16354] = 1'b0;
assign COL[16355] = 1'b0;
assign COL[16356] = 1'b0;
assign COL[16357] = 1'b0;
assign COL[16358] = 1'b0;
assign COL[16359] = 1'b0;
assign COL[16360] = 1'b0;
assign COL[16361] = 1'b0;
assign COL[16362] = 1'b0;
assign COL[16363] = 1'b0;
assign COL[16364] = 1'b0;
assign COL[16365] = 1'b0;
assign COL[16366] = 1'b0;
assign COL[16367] = 1'b0;
assign COL[16368] = 1'b0;
assign COL[16369] = 1'b0;
assign COL[16370] = 1'b0;
assign COL[16371] = 1'b0;
assign COL[16372] = 1'b0;
assign COL[16373] = 1'b0;
assign COL[16374] = 1'b0;
assign COL[16375] = 1'b0;
assign COL[16376] = 1'b0;
assign COL[16377] = 1'b0;
assign COL[16378] = 1'b0;
assign COL[16379] = 1'b0;
assign COL[16380] = 1'b0;
assign COL[16381] = 1'b0;
assign COL[16382] = 1'b0;
assign COL[16383] = 1'b0;
assign COL[16384] = 1'b0;
assign COL[16385] = 1'b0;
assign COL[16386] = 1'b0;
assign COL[16387] = 1'b0;
assign COL[16388] = 1'b0;
assign COL[16389] = 1'b0;
assign COL[16390] = 1'b0;
assign COL[16391] = 1'b0;
assign COL[16392] = 1'b0;
assign COL[16393] = 1'b0;
assign COL[16394] = 1'b0;
assign COL[16395] = 1'b0;
assign COL[16396] = 1'b0;
assign COL[16397] = 1'b0;
assign COL[16398] = 1'b0;
assign COL[16399] = 1'b0;
assign COL[16400] = 1'b0;
assign COL[16401] = 1'b0;
assign COL[16402] = 1'b0;
assign COL[16403] = 1'b0;
assign COL[16404] = 1'b0;
assign COL[16405] = 1'b0;
assign COL[16406] = 1'b0;
assign COL[16407] = 1'b0;
assign COL[16408] = 1'b0;
assign COL[16409] = 1'b0;
assign COL[16410] = 1'b0;
assign COL[16411] = 1'b0;
assign COL[16412] = 1'b0;
assign COL[16413] = 1'b0;
assign COL[16414] = 1'b0;
assign COL[16415] = 1'b0;
assign COL[16416] = 1'b0;
assign COL[16417] = 1'b0;
assign COL[16418] = 1'b0;
assign COL[16419] = 1'b0;
assign COL[16420] = 1'b0;
assign COL[16421] = 1'b0;
assign COL[16422] = 1'b0;
assign COL[16423] = 1'b0;
assign COL[16424] = 1'b0;
assign COL[16425] = 1'b0;
assign COL[16426] = 1'b0;
assign COL[16427] = 1'b0;
assign COL[16428] = 1'b0;
assign COL[16429] = 1'b0;
assign COL[16430] = 1'b0;
assign COL[16431] = 1'b0;
assign COL[16432] = 1'b0;
assign COL[16433] = 1'b0;
assign COL[16434] = 1'b0;
assign COL[16435] = 1'b0;
assign COL[16436] = 1'b0;
assign COL[16437] = 1'b0;
assign COL[16438] = 1'b0;
assign COL[16439] = 1'b0;
assign COL[16440] = 1'b0;
assign COL[16441] = 1'b0;
assign COL[16442] = 1'b0;
assign COL[16443] = 1'b0;
assign COL[16444] = 1'b0;
assign COL[16445] = 1'b0;
assign COL[16446] = 1'b0;
assign COL[16447] = 1'b0;
assign COL[16448] = 1'b0;
assign COL[16449] = 1'b0;
assign COL[16450] = 1'b0;
assign COL[16451] = 1'b0;
assign COL[16452] = 1'b0;
assign COL[16453] = 1'b0;
assign COL[16454] = 1'b0;
assign COL[16455] = 1'b0;
assign COL[16456] = 1'b0;
assign COL[16457] = 1'b0;
assign COL[16458] = 1'b0;
assign COL[16459] = 1'b0;
assign COL[16460] = 1'b0;
assign COL[16461] = 1'b0;
assign COL[16462] = 1'b0;
assign COL[16463] = 1'b0;
assign COL[16464] = 1'b0;
assign COL[16465] = 1'b0;
assign COL[16466] = 1'b0;
assign COL[16467] = 1'b0;
assign COL[16468] = 1'b0;
assign COL[16469] = 1'b0;
assign COL[16470] = 1'b0;
assign COL[16471] = 1'b0;
assign COL[16472] = 1'b0;
assign COL[16473] = 1'b0;
assign COL[16474] = 1'b0;
assign COL[16475] = 1'b0;
assign COL[16476] = 1'b0;
assign COL[16477] = 1'b0;
assign COL[16478] = 1'b0;
assign COL[16479] = 1'b0;
assign COL[16480] = 1'b0;
assign COL[16481] = 1'b0;
assign COL[16482] = 1'b0;
assign COL[16483] = 1'b0;
assign COL[16484] = 1'b0;
assign COL[16485] = 1'b0;
assign COL[16486] = 1'b0;
assign COL[16487] = 1'b0;
assign COL[16488] = 1'b0;
assign COL[16489] = 1'b0;
assign COL[16490] = 1'b0;
assign COL[16491] = 1'b0;
assign COL[16492] = 1'b0;
assign COL[16493] = 1'b0;
assign COL[16494] = 1'b0;
assign COL[16495] = 1'b0;
assign COL[16496] = 1'b0;
assign COL[16497] = 1'b0;
assign COL[16498] = 1'b0;
assign COL[16499] = 1'b0;
assign COL[16500] = 1'b0;
assign COL[16501] = 1'b0;
assign COL[16502] = 1'b0;
assign COL[16503] = 1'b0;
assign COL[16504] = 1'b0;
assign COL[16505] = 1'b0;
assign COL[16506] = 1'b0;
assign COL[16507] = 1'b0;
assign COL[16508] = 1'b0;
assign COL[16509] = 1'b0;
assign COL[16510] = 1'b0;
assign COL[16511] = 1'b0;
assign COL[16512] = 1'b0;
assign COL[16513] = 1'b0;
assign COL[16514] = 1'b0;
assign COL[16515] = 1'b0;
assign COL[16516] = 1'b0;
assign COL[16517] = 1'b0;
assign COL[16518] = 1'b0;
assign COL[16519] = 1'b0;
assign COL[16520] = 1'b0;
assign COL[16521] = 1'b0;
assign COL[16522] = 1'b0;
assign COL[16523] = 1'b0;
assign COL[16524] = 1'b0;
assign COL[16525] = 1'b0;
assign COL[16526] = 1'b0;
assign COL[16527] = 1'b0;
assign COL[16528] = 1'b0;
assign COL[16529] = 1'b0;
assign COL[16530] = 1'b0;
assign COL[16531] = 1'b0;
assign COL[16532] = 1'b0;
assign COL[16533] = 1'b0;
assign COL[16534] = 1'b0;
assign COL[16535] = 1'b0;
assign COL[16536] = 1'b0;
assign COL[16537] = 1'b0;
assign COL[16538] = 1'b0;
assign COL[16539] = 1'b0;
assign COL[16540] = 1'b0;
assign COL[16541] = 1'b0;
assign COL[16542] = 1'b0;
assign COL[16543] = 1'b0;
assign COL[16544] = 1'b0;
assign COL[16545] = 1'b0;
assign COL[16546] = 1'b0;
assign COL[16547] = 1'b0;
assign COL[16548] = 1'b0;
assign COL[16549] = 1'b0;
assign COL[16550] = 1'b0;
assign COL[16551] = 1'b0;
assign COL[16552] = 1'b0;
assign COL[16553] = 1'b0;
assign COL[16554] = 1'b0;
assign COL[16555] = 1'b0;
assign COL[16556] = 1'b0;
assign COL[16557] = 1'b0;
assign COL[16558] = 1'b0;
assign COL[16559] = 1'b0;
assign COL[16560] = 1'b0;
assign COL[16561] = 1'b0;
assign COL[16562] = 1'b0;
assign COL[16563] = 1'b0;
assign COL[16564] = 1'b0;
assign COL[16565] = 1'b0;
assign COL[16566] = 1'b0;
assign COL[16567] = 1'b0;
assign COL[16568] = 1'b0;
assign COL[16569] = 1'b0;
assign COL[16570] = 1'b0;
assign COL[16571] = 1'b0;
assign COL[16572] = 1'b0;
assign COL[16573] = 1'b0;
assign COL[16574] = 1'b0;
assign COL[16575] = 1'b0;
assign COL[16576] = 1'b0;
assign COL[16577] = 1'b0;
assign COL[16578] = 1'b0;
assign COL[16579] = 1'b0;
assign COL[16580] = 1'b0;
assign COL[16581] = 1'b0;
assign COL[16582] = 1'b0;
assign COL[16583] = 1'b0;
assign COL[16584] = 1'b0;
assign COL[16585] = 1'b0;
assign COL[16586] = 1'b0;
assign COL[16587] = 1'b0;
assign COL[16588] = 1'b0;
assign COL[16589] = 1'b0;
assign COL[16590] = 1'b0;
assign COL[16591] = 1'b0;
assign COL[16592] = 1'b0;
assign COL[16593] = 1'b0;
assign COL[16594] = 1'b0;
assign COL[16595] = 1'b0;
assign COL[16596] = 1'b0;
assign COL[16597] = 1'b0;
assign COL[16598] = 1'b0;
assign COL[16599] = 1'b0;
assign COL[16600] = 1'b0;
assign COL[16601] = 1'b0;
assign COL[16602] = 1'b0;
assign COL[16603] = 1'b0;
assign COL[16604] = 1'b0;
assign COL[16605] = 1'b0;
assign COL[16606] = 1'b0;
assign COL[16607] = 1'b0;
assign COL[16608] = 1'b0;
assign COL[16609] = 1'b0;
assign COL[16610] = 1'b0;
assign COL[16611] = 1'b0;
assign COL[16612] = 1'b0;
assign COL[16613] = 1'b0;
assign COL[16614] = 1'b0;
assign COL[16615] = 1'b0;
assign COL[16616] = 1'b0;
assign COL[16617] = 1'b0;
assign COL[16618] = 1'b0;
assign COL[16619] = 1'b0;
assign COL[16620] = 1'b0;
assign COL[16621] = 1'b0;
assign COL[16622] = 1'b0;
assign COL[16623] = 1'b0;
assign COL[16624] = 1'b0;
assign COL[16625] = 1'b0;
assign COL[16626] = 1'b0;
assign COL[16627] = 1'b0;
assign COL[16628] = 1'b0;
assign COL[16629] = 1'b0;
assign COL[16630] = 1'b0;
assign COL[16631] = 1'b0;
assign COL[16632] = 1'b0;
assign COL[16633] = 1'b0;
assign COL[16634] = 1'b0;
assign COL[16635] = 1'b0;
assign COL[16636] = 1'b0;
assign COL[16637] = 1'b0;
assign COL[16638] = 1'b0;
assign COL[16639] = 1'b0;
assign COL[16640] = 1'b0;
assign COL[16641] = 1'b0;
assign COL[16642] = 1'b0;
assign COL[16643] = 1'b0;
assign COL[16644] = 1'b0;
assign COL[16645] = 1'b0;
assign COL[16646] = 1'b0;
assign COL[16647] = 1'b0;
assign COL[16648] = 1'b0;
assign COL[16649] = 1'b0;
assign COL[16650] = 1'b0;
assign COL[16651] = 1'b0;
assign COL[16652] = 1'b0;
assign COL[16653] = 1'b0;
assign COL[16654] = 1'b0;
assign COL[16655] = 1'b0;
assign COL[16656] = 1'b0;
assign COL[16657] = 1'b0;
assign COL[16658] = 1'b0;
assign COL[16659] = 1'b0;
assign COL[16660] = 1'b0;
assign COL[16661] = 1'b0;
assign COL[16662] = 1'b0;
assign COL[16663] = 1'b0;
assign COL[16664] = 1'b0;
assign COL[16665] = 1'b0;
assign COL[16666] = 1'b0;
assign COL[16667] = 1'b0;
assign COL[16668] = 1'b0;
assign COL[16669] = 1'b0;
assign COL[16670] = 1'b0;
assign COL[16671] = 1'b0;
assign COL[16672] = 1'b0;
assign COL[16673] = 1'b0;
assign COL[16674] = 1'b0;
assign COL[16675] = 1'b0;
assign COL[16676] = 1'b0;
assign COL[16677] = 1'b0;
assign COL[16678] = 1'b0;
assign COL[16679] = 1'b0;
assign COL[16680] = 1'b0;
assign COL[16681] = 1'b0;
assign COL[16682] = 1'b0;
assign COL[16683] = 1'b0;
assign COL[16684] = 1'b0;
assign COL[16685] = 1'b0;
assign COL[16686] = 1'b0;
assign COL[16687] = 1'b0;
assign COL[16688] = 1'b0;
assign COL[16689] = 1'b0;
assign COL[16690] = 1'b0;
assign COL[16691] = 1'b0;
assign COL[16692] = 1'b0;
assign COL[16693] = 1'b0;
assign COL[16694] = 1'b0;
assign COL[16695] = 1'b0;
assign COL[16696] = 1'b0;
assign COL[16697] = 1'b0;
assign COL[16698] = 1'b0;
assign COL[16699] = 1'b0;
assign COL[16700] = 1'b0;
assign COL[16701] = 1'b0;
assign COL[16702] = 1'b0;
assign COL[16703] = 1'b0;
assign COL[16704] = 1'b0;
assign COL[16705] = 1'b0;
assign COL[16706] = 1'b0;
assign COL[16707] = 1'b0;
assign COL[16708] = 1'b0;
assign COL[16709] = 1'b0;
assign COL[16710] = 1'b0;
assign COL[16711] = 1'b0;
assign COL[16712] = 1'b0;
assign COL[16713] = 1'b0;
assign COL[16714] = 1'b0;
assign COL[16715] = 1'b0;
assign COL[16716] = 1'b0;
assign COL[16717] = 1'b0;
assign COL[16718] = 1'b0;
assign COL[16719] = 1'b0;
assign COL[16720] = 1'b0;
assign COL[16721] = 1'b0;
assign COL[16722] = 1'b0;
assign COL[16723] = 1'b0;
assign COL[16724] = 1'b0;
assign COL[16725] = 1'b0;
assign COL[16726] = 1'b0;
assign COL[16727] = 1'b0;
assign COL[16728] = 1'b0;
assign COL[16729] = 1'b0;
assign COL[16730] = 1'b0;
assign COL[16731] = 1'b0;
assign COL[16732] = 1'b0;
assign COL[16733] = 1'b0;
assign COL[16734] = 1'b0;
assign COL[16735] = 1'b0;
assign COL[16736] = 1'b0;
assign COL[16737] = 1'b0;
assign COL[16738] = 1'b0;
assign COL[16739] = 1'b0;
assign COL[16740] = 1'b0;
assign COL[16741] = 1'b0;
assign COL[16742] = 1'b0;
assign COL[16743] = 1'b0;
assign COL[16744] = 1'b0;
assign COL[16745] = 1'b0;
assign COL[16746] = 1'b0;
assign COL[16747] = 1'b0;
assign COL[16748] = 1'b0;
assign COL[16749] = 1'b0;
assign COL[16750] = 1'b0;
assign COL[16751] = 1'b0;
assign COL[16752] = 1'b0;
assign COL[16753] = 1'b0;
assign COL[16754] = 1'b0;
assign COL[16755] = 1'b0;
assign COL[16756] = 1'b0;
assign COL[16757] = 1'b0;
assign COL[16758] = 1'b0;
assign COL[16759] = 1'b0;
assign COL[16760] = 1'b0;
assign COL[16761] = 1'b0;
assign COL[16762] = 1'b0;
assign COL[16763] = 1'b0;
assign COL[16764] = 1'b0;
assign COL[16765] = 1'b0;
assign COL[16766] = 1'b0;
assign COL[16767] = 1'b0;
assign COL[16768] = 1'b0;
assign COL[16769] = 1'b0;
assign COL[16770] = 1'b0;
assign COL[16771] = 1'b0;
assign COL[16772] = 1'b0;
assign COL[16773] = 1'b0;
assign COL[16774] = 1'b0;
assign COL[16775] = 1'b0;
assign COL[16776] = 1'b0;
assign COL[16777] = 1'b0;
assign COL[16778] = 1'b0;
assign COL[16779] = 1'b0;
assign COL[16780] = 1'b0;
assign COL[16781] = 1'b0;
assign COL[16782] = 1'b0;
assign COL[16783] = 1'b0;
assign COL[16784] = 1'b0;
assign COL[16785] = 1'b0;
assign COL[16786] = 1'b0;
assign COL[16787] = 1'b0;
assign COL[16788] = 1'b0;
assign COL[16789] = 1'b0;
assign COL[16790] = 1'b0;
assign COL[16791] = 1'b0;
assign COL[16792] = 1'b0;
assign COL[16793] = 1'b0;
assign COL[16794] = 1'b0;
assign COL[16795] = 1'b0;
assign COL[16796] = 1'b0;
assign COL[16797] = 1'b0;
assign COL[16798] = 1'b0;
assign COL[16799] = 1'b0;
assign COL[16800] = 1'b0;
assign COL[16801] = 1'b0;
assign COL[16802] = 1'b0;
assign COL[16803] = 1'b0;
assign COL[16804] = 1'b0;
assign COL[16805] = 1'b0;
assign COL[16806] = 1'b0;
assign COL[16807] = 1'b0;
assign COL[16808] = 1'b0;
assign COL[16809] = 1'b0;
assign COL[16810] = 1'b0;
assign COL[16811] = 1'b0;
assign COL[16812] = 1'b0;
assign COL[16813] = 1'b0;
assign COL[16814] = 1'b0;
assign COL[16815] = 1'b0;
assign COL[16816] = 1'b0;
assign COL[16817] = 1'b0;
assign COL[16818] = 1'b0;
assign COL[16819] = 1'b0;
assign COL[16820] = 1'b0;
assign COL[16821] = 1'b0;
assign COL[16822] = 1'b0;
assign COL[16823] = 1'b0;
assign COL[16824] = 1'b0;
assign COL[16825] = 1'b0;
assign COL[16826] = 1'b0;
assign COL[16827] = 1'b0;
assign COL[16828] = 1'b0;
assign COL[16829] = 1'b0;
assign COL[16830] = 1'b0;
assign COL[16831] = 1'b0;
assign COL[16832] = 1'b0;
assign COL[16833] = 1'b0;
assign COL[16834] = 1'b0;
assign COL[16835] = 1'b0;
assign COL[16836] = 1'b0;
assign COL[16837] = 1'b0;
assign COL[16838] = 1'b0;
assign COL[16839] = 1'b0;
assign COL[16840] = 1'b0;
assign COL[16841] = 1'b0;
assign COL[16842] = 1'b0;
assign COL[16843] = 1'b0;
assign COL[16844] = 1'b0;
assign COL[16845] = 1'b0;
assign COL[16846] = 1'b0;
assign COL[16847] = 1'b0;
assign COL[16848] = 1'b0;
assign COL[16849] = 1'b0;
assign COL[16850] = 1'b0;
assign COL[16851] = 1'b0;
assign COL[16852] = 1'b0;
assign COL[16853] = 1'b0;
assign COL[16854] = 1'b0;
assign COL[16855] = 1'b0;
assign COL[16856] = 1'b0;
assign COL[16857] = 1'b0;
assign COL[16858] = 1'b0;
assign COL[16859] = 1'b0;
assign COL[16860] = 1'b0;
assign COL[16861] = 1'b0;
assign COL[16862] = 1'b0;
assign COL[16863] = 1'b0;
assign COL[16864] = 1'b0;
assign COL[16865] = 1'b0;
assign COL[16866] = 1'b0;
assign COL[16867] = 1'b0;
assign COL[16868] = 1'b0;
assign COL[16869] = 1'b0;
assign COL[16870] = 1'b0;
assign COL[16871] = 1'b0;
assign COL[16872] = 1'b0;
assign COL[16873] = 1'b0;
assign COL[16874] = 1'b0;
assign COL[16875] = 1'b0;
assign COL[16876] = 1'b0;
assign COL[16877] = 1'b0;
assign COL[16878] = 1'b0;
assign COL[16879] = 1'b0;
assign COL[16880] = 1'b0;
assign COL[16881] = 1'b0;
assign COL[16882] = 1'b0;
assign COL[16883] = 1'b0;
assign COL[16884] = 1'b0;
assign COL[16885] = 1'b0;
assign COL[16886] = 1'b0;
assign COL[16887] = 1'b0;
assign COL[16888] = 1'b0;
assign COL[16889] = 1'b0;
assign COL[16890] = 1'b0;
assign COL[16891] = 1'b0;
assign COL[16892] = 1'b0;
assign COL[16893] = 1'b0;
assign COL[16894] = 1'b0;
assign COL[16895] = 1'b0;
assign COL[16896] = 1'b0;
assign COL[16897] = 1'b0;
assign COL[16898] = 1'b0;
assign COL[16899] = 1'b0;
assign COL[16900] = 1'b0;
assign COL[16901] = 1'b0;
assign COL[16902] = 1'b0;
assign COL[16903] = 1'b0;
assign COL[16904] = 1'b0;
assign COL[16905] = 1'b0;
assign COL[16906] = 1'b0;
assign COL[16907] = 1'b0;
assign COL[16908] = 1'b0;
assign COL[16909] = 1'b0;
assign COL[16910] = 1'b0;
assign COL[16911] = 1'b0;
assign COL[16912] = 1'b0;
assign COL[16913] = 1'b0;
assign COL[16914] = 1'b0;
assign COL[16915] = 1'b0;
assign COL[16916] = 1'b0;
assign COL[16917] = 1'b0;
assign COL[16918] = 1'b0;
assign COL[16919] = 1'b0;
assign COL[16920] = 1'b0;
assign COL[16921] = 1'b0;
assign COL[16922] = 1'b0;
assign COL[16923] = 1'b0;
assign COL[16924] = 1'b0;
assign COL[16925] = 1'b0;
assign COL[16926] = 1'b0;
assign COL[16927] = 1'b0;
assign COL[16928] = 1'b0;
assign COL[16929] = 1'b0;
assign COL[16930] = 1'b0;
assign COL[16931] = 1'b0;
assign COL[16932] = 1'b0;
assign COL[16933] = 1'b0;
assign COL[16934] = 1'b0;
assign COL[16935] = 1'b0;
assign COL[16936] = 1'b0;
assign COL[16937] = 1'b0;
assign COL[16938] = 1'b0;
assign COL[16939] = 1'b0;
assign COL[16940] = 1'b0;
assign COL[16941] = 1'b0;
assign COL[16942] = 1'b0;
assign COL[16943] = 1'b0;
assign COL[16944] = 1'b0;
assign COL[16945] = 1'b0;
assign COL[16946] = 1'b0;
assign COL[16947] = 1'b0;
assign COL[16948] = 1'b0;
assign COL[16949] = 1'b0;
assign COL[16950] = 1'b0;
assign COL[16951] = 1'b0;
assign COL[16952] = 1'b0;
assign COL[16953] = 1'b0;
assign COL[16954] = 1'b0;
assign COL[16955] = 1'b0;
assign COL[16956] = 1'b0;
assign COL[16957] = 1'b0;
assign COL[16958] = 1'b0;
assign COL[16959] = 1'b0;
assign COL[16960] = 1'b0;
assign COL[16961] = 1'b0;
assign COL[16962] = 1'b0;
assign COL[16963] = 1'b0;
assign COL[16964] = 1'b0;
assign COL[16965] = 1'b0;
assign COL[16966] = 1'b0;
assign COL[16967] = 1'b0;
assign COL[16968] = 1'b0;
assign COL[16969] = 1'b0;
assign COL[16970] = 1'b0;
assign COL[16971] = 1'b0;
assign COL[16972] = 1'b0;
assign COL[16973] = 1'b0;
assign COL[16974] = 1'b0;
assign COL[16975] = 1'b0;
assign COL[16976] = 1'b0;
assign COL[16977] = 1'b0;
assign COL[16978] = 1'b0;
assign COL[16979] = 1'b0;
assign COL[16980] = 1'b0;
assign COL[16981] = 1'b0;
assign COL[16982] = 1'b0;
assign COL[16983] = 1'b0;
assign COL[16984] = 1'b0;
assign COL[16985] = 1'b0;
assign COL[16986] = 1'b0;
assign COL[16987] = 1'b0;
assign COL[16988] = 1'b0;
assign COL[16989] = 1'b0;
assign COL[16990] = 1'b0;
assign COL[16991] = 1'b0;
assign COL[16992] = 1'b0;
assign COL[16993] = 1'b0;
assign COL[16994] = 1'b0;
assign COL[16995] = 1'b0;
assign COL[16996] = 1'b0;
assign COL[16997] = 1'b0;
assign COL[16998] = 1'b0;
assign COL[16999] = 1'b0;
assign COL[17000] = 1'b0;
assign COL[17001] = 1'b0;
assign COL[17002] = 1'b0;
assign COL[17003] = 1'b0;
assign COL[17004] = 1'b0;
assign COL[17005] = 1'b0;
assign COL[17006] = 1'b0;
assign COL[17007] = 1'b0;
assign COL[17008] = 1'b0;
assign COL[17009] = 1'b0;
assign COL[17010] = 1'b0;
assign COL[17011] = 1'b0;
assign COL[17012] = 1'b0;
assign COL[17013] = 1'b0;
assign COL[17014] = 1'b0;
assign COL[17015] = 1'b0;
assign COL[17016] = 1'b0;
assign COL[17017] = 1'b0;
assign COL[17018] = 1'b0;
assign COL[17019] = 1'b0;
assign COL[17020] = 1'b0;
assign COL[17021] = 1'b0;
assign COL[17022] = 1'b0;
assign COL[17023] = 1'b0;
assign COL[17024] = 1'b0;
assign COL[17025] = 1'b0;
assign COL[17026] = 1'b0;
assign COL[17027] = 1'b0;
assign COL[17028] = 1'b0;
assign COL[17029] = 1'b0;
assign COL[17030] = 1'b0;
assign COL[17031] = 1'b0;
assign COL[17032] = 1'b0;
assign COL[17033] = 1'b0;
assign COL[17034] = 1'b0;
assign COL[17035] = 1'b0;
assign COL[17036] = 1'b0;
assign COL[17037] = 1'b0;
assign COL[17038] = 1'b0;
assign COL[17039] = 1'b0;
assign COL[17040] = 1'b0;
assign COL[17041] = 1'b0;
assign COL[17042] = 1'b0;
assign COL[17043] = 1'b0;
assign COL[17044] = 1'b0;
assign COL[17045] = 1'b0;
assign COL[17046] = 1'b0;
assign COL[17047] = 1'b0;
assign COL[17048] = 1'b0;
assign COL[17049] = 1'b0;
assign COL[17050] = 1'b0;
assign COL[17051] = 1'b0;
assign COL[17052] = 1'b0;
assign COL[17053] = 1'b0;
assign COL[17054] = 1'b0;
assign COL[17055] = 1'b0;
assign COL[17056] = 1'b0;
assign COL[17057] = 1'b0;
assign COL[17058] = 1'b0;
assign COL[17059] = 1'b0;
assign COL[17060] = 1'b0;
assign COL[17061] = 1'b0;
assign COL[17062] = 1'b0;
assign COL[17063] = 1'b0;
assign COL[17064] = 1'b0;
assign COL[17065] = 1'b0;
assign COL[17066] = 1'b0;
assign COL[17067] = 1'b0;
assign COL[17068] = 1'b0;
assign COL[17069] = 1'b0;
assign COL[17070] = 1'b0;
assign COL[17071] = 1'b0;
assign COL[17072] = 1'b0;
assign COL[17073] = 1'b0;
assign COL[17074] = 1'b0;
assign COL[17075] = 1'b0;
assign COL[17076] = 1'b0;
assign COL[17077] = 1'b0;
assign COL[17078] = 1'b0;
assign COL[17079] = 1'b0;
assign COL[17080] = 1'b0;
assign COL[17081] = 1'b0;
assign COL[17082] = 1'b0;
assign COL[17083] = 1'b0;
assign COL[17084] = 1'b0;
assign COL[17085] = 1'b0;
assign COL[17086] = 1'b0;
assign COL[17087] = 1'b0;
assign COL[17088] = 1'b0;
assign COL[17089] = 1'b0;
assign COL[17090] = 1'b0;
assign COL[17091] = 1'b0;
assign COL[17092] = 1'b0;
assign COL[17093] = 1'b0;
assign COL[17094] = 1'b0;
assign COL[17095] = 1'b0;
assign COL[17096] = 1'b0;
assign COL[17097] = 1'b0;
assign COL[17098] = 1'b0;
assign COL[17099] = 1'b0;
assign COL[17100] = 1'b0;
assign COL[17101] = 1'b0;
assign COL[17102] = 1'b0;
assign COL[17103] = 1'b0;
assign COL[17104] = 1'b0;
assign COL[17105] = 1'b0;
assign COL[17106] = 1'b0;
assign COL[17107] = 1'b0;
assign COL[17108] = 1'b0;
assign COL[17109] = 1'b0;
assign COL[17110] = 1'b0;
assign COL[17111] = 1'b0;
assign COL[17112] = 1'b0;
assign COL[17113] = 1'b0;
assign COL[17114] = 1'b0;
assign COL[17115] = 1'b0;
assign COL[17116] = 1'b0;
assign COL[17117] = 1'b0;
assign COL[17118] = 1'b0;
assign COL[17119] = 1'b0;
assign COL[17120] = 1'b0;
assign COL[17121] = 1'b0;
assign COL[17122] = 1'b0;
assign COL[17123] = 1'b0;
assign COL[17124] = 1'b0;
assign COL[17125] = 1'b0;
assign COL[17126] = 1'b0;
assign COL[17127] = 1'b0;
assign COL[17128] = 1'b0;
assign COL[17129] = 1'b0;
assign COL[17130] = 1'b0;
assign COL[17131] = 1'b0;
assign COL[17132] = 1'b0;
assign COL[17133] = 1'b0;
assign COL[17134] = 1'b0;
assign COL[17135] = 1'b0;
assign COL[17136] = 1'b0;
assign COL[17137] = 1'b0;
assign COL[17138] = 1'b0;
assign COL[17139] = 1'b0;
assign COL[17140] = 1'b0;
assign COL[17141] = 1'b0;
assign COL[17142] = 1'b0;
assign COL[17143] = 1'b0;
assign COL[17144] = 1'b0;
assign COL[17145] = 1'b0;
assign COL[17146] = 1'b0;
assign COL[17147] = 1'b0;
assign COL[17148] = 1'b0;
assign COL[17149] = 1'b0;
assign COL[17150] = 1'b0;
assign COL[17151] = 1'b0;
assign COL[17152] = 1'b0;
assign COL[17153] = 1'b0;
assign COL[17154] = 1'b0;
assign COL[17155] = 1'b0;
assign COL[17156] = 1'b0;
assign COL[17157] = 1'b0;
assign COL[17158] = 1'b0;
assign COL[17159] = 1'b0;
assign COL[17160] = 1'b0;
assign COL[17161] = 1'b0;
assign COL[17162] = 1'b0;
assign COL[17163] = 1'b0;
assign COL[17164] = 1'b0;
assign COL[17165] = 1'b0;
assign COL[17166] = 1'b0;
assign COL[17167] = 1'b0;
assign COL[17168] = 1'b0;
assign COL[17169] = 1'b0;
assign COL[17170] = 1'b0;
assign COL[17171] = 1'b0;
assign COL[17172] = 1'b0;
assign COL[17173] = 1'b0;
assign COL[17174] = 1'b0;
assign COL[17175] = 1'b0;
assign COL[17176] = 1'b0;
assign COL[17177] = 1'b0;
assign COL[17178] = 1'b0;
assign COL[17179] = 1'b0;
assign COL[17180] = 1'b0;
assign COL[17181] = 1'b0;
assign COL[17182] = 1'b0;
assign COL[17183] = 1'b0;
assign COL[17184] = 1'b0;
assign COL[17185] = 1'b0;
assign COL[17186] = 1'b0;
assign COL[17187] = 1'b0;
assign COL[17188] = 1'b0;
assign COL[17189] = 1'b0;
assign COL[17190] = 1'b0;
assign COL[17191] = 1'b0;
assign COL[17192] = 1'b0;
assign COL[17193] = 1'b0;
assign COL[17194] = 1'b0;
assign COL[17195] = 1'b0;
assign COL[17196] = 1'b0;
assign COL[17197] = 1'b0;
assign COL[17198] = 1'b0;
assign COL[17199] = 1'b0;
assign COL[17200] = 1'b0;
assign COL[17201] = 1'b0;
assign COL[17202] = 1'b0;
assign COL[17203] = 1'b0;
assign COL[17204] = 1'b0;
assign COL[17205] = 1'b0;
assign COL[17206] = 1'b0;
assign COL[17207] = 1'b0;
assign COL[17208] = 1'b0;
assign COL[17209] = 1'b0;
assign COL[17210] = 1'b0;
assign COL[17211] = 1'b0;
assign COL[17212] = 1'b0;
assign COL[17213] = 1'b0;
assign COL[17214] = 1'b0;
assign COL[17215] = 1'b0;
assign COL[17216] = 1'b0;
assign COL[17217] = 1'b0;
assign COL[17218] = 1'b0;
assign COL[17219] = 1'b0;
assign COL[17220] = 1'b0;
assign COL[17221] = 1'b0;
assign COL[17222] = 1'b0;
assign COL[17223] = 1'b0;
assign COL[17224] = 1'b0;
assign COL[17225] = 1'b0;
assign COL[17226] = 1'b0;
assign COL[17227] = 1'b0;
assign COL[17228] = 1'b0;
assign COL[17229] = 1'b0;
assign COL[17230] = 1'b0;
assign COL[17231] = 1'b0;
assign COL[17232] = 1'b0;
assign COL[17233] = 1'b0;
assign COL[17234] = 1'b0;
assign COL[17235] = 1'b0;
assign COL[17236] = 1'b0;
assign COL[17237] = 1'b0;
assign COL[17238] = 1'b0;
assign COL[17239] = 1'b0;
assign COL[17240] = 1'b0;
assign COL[17241] = 1'b0;
assign COL[17242] = 1'b0;
assign COL[17243] = 1'b0;
assign COL[17244] = 1'b0;
assign COL[17245] = 1'b0;
assign COL[17246] = 1'b0;
assign COL[17247] = 1'b0;
assign COL[17248] = 1'b0;
assign COL[17249] = 1'b0;
assign COL[17250] = 1'b0;
assign COL[17251] = 1'b0;
assign COL[17252] = 1'b0;
assign COL[17253] = 1'b0;
assign COL[17254] = 1'b0;
assign COL[17255] = 1'b0;
assign COL[17256] = 1'b0;
assign COL[17257] = 1'b0;
assign COL[17258] = 1'b0;
assign COL[17259] = 1'b0;
assign COL[17260] = 1'b0;
assign COL[17261] = 1'b0;
assign COL[17262] = 1'b0;
assign COL[17263] = 1'b0;
assign COL[17264] = 1'b0;
assign COL[17265] = 1'b0;
assign COL[17266] = 1'b0;
assign COL[17267] = 1'b0;
assign COL[17268] = 1'b0;
assign COL[17269] = 1'b0;
assign COL[17270] = 1'b0;
assign COL[17271] = 1'b0;
assign COL[17272] = 1'b0;
assign COL[17273] = 1'b0;
assign COL[17274] = 1'b0;
assign COL[17275] = 1'b0;
assign COL[17276] = 1'b0;
assign COL[17277] = 1'b0;
assign COL[17278] = 1'b0;
assign COL[17279] = 1'b0;
assign COL[17280] = 1'b0;
assign COL[17281] = 1'b0;
assign COL[17282] = 1'b0;
assign COL[17283] = 1'b0;
assign COL[17284] = 1'b0;
assign COL[17285] = 1'b0;
assign COL[17286] = 1'b0;
assign COL[17287] = 1'b0;
assign COL[17288] = 1'b0;
assign COL[17289] = 1'b0;
assign COL[17290] = 1'b0;
assign COL[17291] = 1'b0;
assign COL[17292] = 1'b0;
assign COL[17293] = 1'b0;
assign COL[17294] = 1'b0;
assign COL[17295] = 1'b0;
assign COL[17296] = 1'b0;
assign COL[17297] = 1'b0;
assign COL[17298] = 1'b0;
assign COL[17299] = 1'b0;
assign COL[17300] = 1'b0;
assign COL[17301] = 1'b0;
assign COL[17302] = 1'b0;
assign COL[17303] = 1'b0;
assign COL[17304] = 1'b0;
assign COL[17305] = 1'b0;
assign COL[17306] = 1'b0;
assign COL[17307] = 1'b0;
assign COL[17308] = 1'b0;
assign COL[17309] = 1'b0;
assign COL[17310] = 1'b0;
assign COL[17311] = 1'b0;
assign COL[17312] = 1'b0;
assign COL[17313] = 1'b0;
assign COL[17314] = 1'b0;
assign COL[17315] = 1'b0;
assign COL[17316] = 1'b0;
assign COL[17317] = 1'b0;
assign COL[17318] = 1'b0;
assign COL[17319] = 1'b0;
assign COL[17320] = 1'b0;
assign COL[17321] = 1'b0;
assign COL[17322] = 1'b0;
assign COL[17323] = 1'b0;
assign COL[17324] = 1'b0;
assign COL[17325] = 1'b0;
assign COL[17326] = 1'b0;
assign COL[17327] = 1'b0;
assign COL[17328] = 1'b0;
assign COL[17329] = 1'b0;
assign COL[17330] = 1'b0;
assign COL[17331] = 1'b0;
assign COL[17332] = 1'b0;
assign COL[17333] = 1'b0;
assign COL[17334] = 1'b0;
assign COL[17335] = 1'b0;
assign COL[17336] = 1'b0;
assign COL[17337] = 1'b0;
assign COL[17338] = 1'b0;
assign COL[17339] = 1'b0;
assign COL[17340] = 1'b0;
assign COL[17341] = 1'b0;
assign COL[17342] = 1'b0;
assign COL[17343] = 1'b0;
assign COL[17344] = 1'b0;
assign COL[17345] = 1'b0;
assign COL[17346] = 1'b0;
assign COL[17347] = 1'b0;
assign COL[17348] = 1'b0;
assign COL[17349] = 1'b0;
assign COL[17350] = 1'b0;
assign COL[17351] = 1'b0;
assign COL[17352] = 1'b0;
assign COL[17353] = 1'b0;
assign COL[17354] = 1'b0;
assign COL[17355] = 1'b0;
assign COL[17356] = 1'b0;
assign COL[17357] = 1'b0;
assign COL[17358] = 1'b0;
assign COL[17359] = 1'b0;
assign COL[17360] = 1'b0;
assign COL[17361] = 1'b0;
assign COL[17362] = 1'b0;
assign COL[17363] = 1'b0;
assign COL[17364] = 1'b0;
assign COL[17365] = 1'b0;
assign COL[17366] = 1'b0;
assign COL[17367] = 1'b0;
assign COL[17368] = 1'b0;
assign COL[17369] = 1'b0;
assign COL[17370] = 1'b0;
assign COL[17371] = 1'b0;
assign COL[17372] = 1'b0;
assign COL[17373] = 1'b0;
assign COL[17374] = 1'b0;
assign COL[17375] = 1'b0;
assign COL[17376] = 1'b0;
assign COL[17377] = 1'b0;
assign COL[17378] = 1'b0;
assign COL[17379] = 1'b0;
assign COL[17380] = 1'b0;
assign COL[17381] = 1'b0;
assign COL[17382] = 1'b0;
assign COL[17383] = 1'b0;
assign COL[17384] = 1'b0;
assign COL[17385] = 1'b0;
assign COL[17386] = 1'b0;
assign COL[17387] = 1'b0;
assign COL[17388] = 1'b0;
assign COL[17389] = 1'b0;
assign COL[17390] = 1'b0;
assign COL[17391] = 1'b0;
assign COL[17392] = 1'b0;
assign COL[17393] = 1'b0;
assign COL[17394] = 1'b0;
assign COL[17395] = 1'b0;
assign COL[17396] = 1'b0;
assign COL[17397] = 1'b0;
assign COL[17398] = 1'b0;
assign COL[17399] = 1'b0;
assign COL[17400] = 1'b0;
assign COL[17401] = 1'b0;
assign COL[17402] = 1'b0;
assign COL[17403] = 1'b0;
assign COL[17404] = 1'b0;
assign COL[17405] = 1'b0;
assign COL[17406] = 1'b0;
assign COL[17407] = 1'b0;
assign COL[17408] = 1'b0;
assign COL[17409] = 1'b0;
assign COL[17410] = 1'b0;
assign COL[17411] = 1'b0;
assign COL[17412] = 1'b0;
assign COL[17413] = 1'b0;
assign COL[17414] = 1'b0;
assign COL[17415] = 1'b0;
assign COL[17416] = 1'b0;
assign COL[17417] = 1'b0;
assign COL[17418] = 1'b0;
assign COL[17419] = 1'b0;
assign COL[17420] = 1'b0;
assign COL[17421] = 1'b0;
assign COL[17422] = 1'b0;
assign COL[17423] = 1'b0;
assign COL[17424] = 1'b0;
assign COL[17425] = 1'b0;
assign COL[17426] = 1'b0;
assign COL[17427] = 1'b0;
assign COL[17428] = 1'b0;
assign COL[17429] = 1'b0;
assign COL[17430] = 1'b0;
assign COL[17431] = 1'b0;
assign COL[17432] = 1'b0;
assign COL[17433] = 1'b0;
assign COL[17434] = 1'b0;
assign COL[17435] = 1'b0;
assign COL[17436] = 1'b0;
assign COL[17437] = 1'b0;
assign COL[17438] = 1'b0;
assign COL[17439] = 1'b0;
assign COL[17440] = 1'b0;
assign COL[17441] = 1'b0;
assign COL[17442] = 1'b0;
assign COL[17443] = 1'b0;
assign COL[17444] = 1'b0;
assign COL[17445] = 1'b0;
assign COL[17446] = 1'b0;
assign COL[17447] = 1'b0;
assign COL[17448] = 1'b0;
assign COL[17449] = 1'b0;
assign COL[17450] = 1'b0;
assign COL[17451] = 1'b0;
assign COL[17452] = 1'b0;
assign COL[17453] = 1'b0;
assign COL[17454] = 1'b0;
assign COL[17455] = 1'b0;
assign COL[17456] = 1'b0;
assign COL[17457] = 1'b0;
assign COL[17458] = 1'b0;
assign COL[17459] = 1'b0;
assign COL[17460] = 1'b0;
assign COL[17461] = 1'b0;
assign COL[17462] = 1'b0;
assign COL[17463] = 1'b0;
assign COL[17464] = 1'b0;
assign COL[17465] = 1'b0;
assign COL[17466] = 1'b0;
assign COL[17467] = 1'b0;
assign COL[17468] = 1'b0;
assign COL[17469] = 1'b0;
assign COL[17470] = 1'b0;
assign COL[17471] = 1'b0;
assign COL[17472] = 1'b0;
assign COL[17473] = 1'b0;
assign COL[17474] = 1'b0;
assign COL[17475] = 1'b0;
assign COL[17476] = 1'b0;
assign COL[17477] = 1'b0;
assign COL[17478] = 1'b0;
assign COL[17479] = 1'b0;
assign COL[17480] = 1'b0;
assign COL[17481] = 1'b0;
assign COL[17482] = 1'b0;
assign COL[17483] = 1'b0;
assign COL[17484] = 1'b0;
assign COL[17485] = 1'b0;
assign COL[17486] = 1'b0;
assign COL[17487] = 1'b0;
assign COL[17488] = 1'b0;
assign COL[17489] = 1'b0;
assign COL[17490] = 1'b0;
assign COL[17491] = 1'b0;
assign COL[17492] = 1'b0;
assign COL[17493] = 1'b0;
assign COL[17494] = 1'b0;
assign COL[17495] = 1'b0;
assign COL[17496] = 1'b0;
assign COL[17497] = 1'b0;
assign COL[17498] = 1'b0;
assign COL[17499] = 1'b0;
assign COL[17500] = 1'b0;
assign COL[17501] = 1'b0;
assign COL[17502] = 1'b0;
assign COL[17503] = 1'b0;
assign COL[17504] = 1'b0;
assign COL[17505] = 1'b0;
assign COL[17506] = 1'b0;
assign COL[17507] = 1'b0;
assign COL[17508] = 1'b0;
assign COL[17509] = 1'b0;
assign COL[17510] = 1'b0;
assign COL[17511] = 1'b0;
assign COL[17512] = 1'b0;
assign COL[17513] = 1'b0;
assign COL[17514] = 1'b0;
assign COL[17515] = 1'b0;
assign COL[17516] = 1'b0;
assign COL[17517] = 1'b0;
assign COL[17518] = 1'b0;
assign COL[17519] = 1'b0;
assign COL[17520] = 1'b0;
assign COL[17521] = 1'b0;
assign COL[17522] = 1'b0;
assign COL[17523] = 1'b0;
assign COL[17524] = 1'b0;
assign COL[17525] = 1'b0;
assign COL[17526] = 1'b0;
assign COL[17527] = 1'b0;
assign COL[17528] = 1'b0;
assign COL[17529] = 1'b0;
assign COL[17530] = 1'b0;
assign COL[17531] = 1'b0;
assign COL[17532] = 1'b0;
assign COL[17533] = 1'b0;
assign COL[17534] = 1'b0;
assign COL[17535] = 1'b0;
assign COL[17536] = 1'b0;
assign COL[17537] = 1'b0;
assign COL[17538] = 1'b0;
assign COL[17539] = 1'b0;
assign COL[17540] = 1'b0;
assign COL[17541] = 1'b0;
assign COL[17542] = 1'b0;
assign COL[17543] = 1'b0;
assign COL[17544] = 1'b0;
assign COL[17545] = 1'b0;
assign COL[17546] = 1'b0;
assign COL[17547] = 1'b0;
assign COL[17548] = 1'b0;
assign COL[17549] = 1'b0;
assign COL[17550] = 1'b0;
assign COL[17551] = 1'b0;
assign COL[17552] = 1'b0;
assign COL[17553] = 1'b0;
assign COL[17554] = 1'b0;
assign COL[17555] = 1'b0;
assign COL[17556] = 1'b0;
assign COL[17557] = 1'b0;
assign COL[17558] = 1'b0;
assign COL[17559] = 1'b0;
assign COL[17560] = 1'b0;
assign COL[17561] = 1'b0;
assign COL[17562] = 1'b0;
assign COL[17563] = 1'b0;
assign COL[17564] = 1'b0;
assign COL[17565] = 1'b0;
assign COL[17566] = 1'b0;
assign COL[17567] = 1'b0;
assign COL[17568] = 1'b0;
assign COL[17569] = 1'b0;
assign COL[17570] = 1'b0;
assign COL[17571] = 1'b0;
assign COL[17572] = 1'b0;
assign COL[17573] = 1'b0;
assign COL[17574] = 1'b0;
assign COL[17575] = 1'b0;
assign COL[17576] = 1'b0;
assign COL[17577] = 1'b0;
assign COL[17578] = 1'b0;
assign COL[17579] = 1'b0;
assign COL[17580] = 1'b0;
assign COL[17581] = 1'b0;
assign COL[17582] = 1'b0;
assign COL[17583] = 1'b0;
assign COL[17584] = 1'b0;
assign COL[17585] = 1'b0;
assign COL[17586] = 1'b0;
assign COL[17587] = 1'b0;
assign COL[17588] = 1'b0;
assign COL[17589] = 1'b0;
assign COL[17590] = 1'b0;
assign COL[17591] = 1'b0;
assign COL[17592] = 1'b0;
assign COL[17593] = 1'b0;
assign COL[17594] = 1'b0;
assign COL[17595] = 1'b0;
assign COL[17596] = 1'b0;
assign COL[17597] = 1'b0;
assign COL[17598] = 1'b0;
assign COL[17599] = 1'b0;
assign COL[17600] = 1'b0;
assign COL[17601] = 1'b0;
assign COL[17602] = 1'b0;
assign COL[17603] = 1'b0;
assign COL[17604] = 1'b0;
assign COL[17605] = 1'b0;
assign COL[17606] = 1'b0;
assign COL[17607] = 1'b0;
assign COL[17608] = 1'b0;
assign COL[17609] = 1'b0;
assign COL[17610] = 1'b0;
assign COL[17611] = 1'b0;
assign COL[17612] = 1'b0;
assign COL[17613] = 1'b0;
assign COL[17614] = 1'b0;
assign COL[17615] = 1'b0;
assign COL[17616] = 1'b0;
assign COL[17617] = 1'b0;
assign COL[17618] = 1'b0;
assign COL[17619] = 1'b0;
assign COL[17620] = 1'b0;
assign COL[17621] = 1'b0;
assign COL[17622] = 1'b0;
assign COL[17623] = 1'b0;
assign COL[17624] = 1'b0;
assign COL[17625] = 1'b0;
assign COL[17626] = 1'b0;
assign COL[17627] = 1'b0;
assign COL[17628] = 1'b0;
assign COL[17629] = 1'b0;
assign COL[17630] = 1'b0;
assign COL[17631] = 1'b0;
assign COL[17632] = 1'b0;
assign COL[17633] = 1'b0;
assign COL[17634] = 1'b0;
assign COL[17635] = 1'b0;
assign COL[17636] = 1'b0;
assign COL[17637] = 1'b0;
assign COL[17638] = 1'b0;
assign COL[17639] = 1'b0;
assign COL[17640] = 1'b0;
assign COL[17641] = 1'b0;
assign COL[17642] = 1'b0;
assign COL[17643] = 1'b0;
assign COL[17644] = 1'b0;
assign COL[17645] = 1'b0;
assign COL[17646] = 1'b0;
assign COL[17647] = 1'b0;
assign COL[17648] = 1'b0;
assign COL[17649] = 1'b0;
assign COL[17650] = 1'b0;
assign COL[17651] = 1'b0;
assign COL[17652] = 1'b0;
assign COL[17653] = 1'b0;
assign COL[17654] = 1'b0;
assign COL[17655] = 1'b0;
assign COL[17656] = 1'b0;
assign COL[17657] = 1'b0;
assign COL[17658] = 1'b0;
assign COL[17659] = 1'b0;
assign COL[17660] = 1'b0;
assign COL[17661] = 1'b0;
assign COL[17662] = 1'b0;
assign COL[17663] = 1'b0;
assign COL[17664] = 1'b0;
assign COL[17665] = 1'b0;
assign COL[17666] = 1'b0;
assign COL[17667] = 1'b0;
assign COL[17668] = 1'b0;
assign COL[17669] = 1'b0;
assign COL[17670] = 1'b0;
assign COL[17671] = 1'b0;
assign COL[17672] = 1'b0;
assign COL[17673] = 1'b0;
assign COL[17674] = 1'b0;
assign COL[17675] = 1'b0;
assign COL[17676] = 1'b0;
assign COL[17677] = 1'b0;
assign COL[17678] = 1'b0;
assign COL[17679] = 1'b0;
assign COL[17680] = 1'b0;
assign COL[17681] = 1'b0;
assign COL[17682] = 1'b0;
assign COL[17683] = 1'b0;
assign COL[17684] = 1'b0;
assign COL[17685] = 1'b0;
assign COL[17686] = 1'b0;
assign COL[17687] = 1'b0;
assign COL[17688] = 1'b0;
assign COL[17689] = 1'b0;
assign COL[17690] = 1'b0;
assign COL[17691] = 1'b0;
assign COL[17692] = 1'b0;
assign COL[17693] = 1'b0;
assign COL[17694] = 1'b0;
assign COL[17695] = 1'b0;
assign COL[17696] = 1'b0;
assign COL[17697] = 1'b0;
assign COL[17698] = 1'b0;
assign COL[17699] = 1'b0;
assign COL[17700] = 1'b0;
assign COL[17701] = 1'b0;
assign COL[17702] = 1'b0;
assign COL[17703] = 1'b0;
assign COL[17704] = 1'b0;
assign COL[17705] = 1'b0;
assign COL[17706] = 1'b0;
assign COL[17707] = 1'b0;
assign COL[17708] = 1'b0;
assign COL[17709] = 1'b0;
assign COL[17710] = 1'b0;
assign COL[17711] = 1'b0;
assign COL[17712] = 1'b0;
assign COL[17713] = 1'b0;
assign COL[17714] = 1'b0;
assign COL[17715] = 1'b0;
assign COL[17716] = 1'b0;
assign COL[17717] = 1'b0;
assign COL[17718] = 1'b0;
assign COL[17719] = 1'b0;
assign COL[17720] = 1'b0;
assign COL[17721] = 1'b0;
assign COL[17722] = 1'b0;
assign COL[17723] = 1'b0;
assign COL[17724] = 1'b0;
assign COL[17725] = 1'b0;
assign COL[17726] = 1'b0;
assign COL[17727] = 1'b0;
assign COL[17728] = 1'b0;
assign COL[17729] = 1'b0;
assign COL[17730] = 1'b0;
assign COL[17731] = 1'b0;
assign COL[17732] = 1'b0;
assign COL[17733] = 1'b0;
assign COL[17734] = 1'b0;
assign COL[17735] = 1'b0;
assign COL[17736] = 1'b0;
assign COL[17737] = 1'b0;
assign COL[17738] = 1'b0;
assign COL[17739] = 1'b0;
assign COL[17740] = 1'b0;
assign COL[17741] = 1'b0;
assign COL[17742] = 1'b0;
assign COL[17743] = 1'b0;
assign COL[17744] = 1'b0;
assign COL[17745] = 1'b0;
assign COL[17746] = 1'b0;
assign COL[17747] = 1'b0;
assign COL[17748] = 1'b0;
assign COL[17749] = 1'b0;
assign COL[17750] = 1'b0;
assign COL[17751] = 1'b0;
assign COL[17752] = 1'b0;
assign COL[17753] = 1'b0;
assign COL[17754] = 1'b0;
assign COL[17755] = 1'b0;
assign COL[17756] = 1'b0;
assign COL[17757] = 1'b0;
assign COL[17758] = 1'b0;
assign COL[17759] = 1'b0;
assign COL[17760] = 1'b0;
assign COL[17761] = 1'b0;
assign COL[17762] = 1'b0;
assign COL[17763] = 1'b0;
assign COL[17764] = 1'b0;
assign COL[17765] = 1'b0;
assign COL[17766] = 1'b0;
assign COL[17767] = 1'b0;
assign COL[17768] = 1'b0;
assign COL[17769] = 1'b0;
assign COL[17770] = 1'b0;
assign COL[17771] = 1'b0;
assign COL[17772] = 1'b0;
assign COL[17773] = 1'b0;
assign COL[17774] = 1'b0;
assign COL[17775] = 1'b0;
assign COL[17776] = 1'b0;
assign COL[17777] = 1'b0;
assign COL[17778] = 1'b0;
assign COL[17779] = 1'b0;
assign COL[17780] = 1'b0;
assign COL[17781] = 1'b0;
assign COL[17782] = 1'b0;
assign COL[17783] = 1'b0;
assign COL[17784] = 1'b0;
assign COL[17785] = 1'b0;
assign COL[17786] = 1'b0;
assign COL[17787] = 1'b0;
assign COL[17788] = 1'b0;
assign COL[17789] = 1'b0;
assign COL[17790] = 1'b0;
assign COL[17791] = 1'b0;
assign COL[17792] = 1'b0;
assign COL[17793] = 1'b0;
assign COL[17794] = 1'b0;
assign COL[17795] = 1'b0;
assign COL[17796] = 1'b0;
assign COL[17797] = 1'b0;
assign COL[17798] = 1'b0;
assign COL[17799] = 1'b0;
assign COL[17800] = 1'b0;
assign COL[17801] = 1'b0;
assign COL[17802] = 1'b0;
assign COL[17803] = 1'b0;
assign COL[17804] = 1'b0;
assign COL[17805] = 1'b0;
assign COL[17806] = 1'b0;
assign COL[17807] = 1'b0;
assign COL[17808] = 1'b0;
assign COL[17809] = 1'b0;
assign COL[17810] = 1'b0;
assign COL[17811] = 1'b0;
assign COL[17812] = 1'b0;
assign COL[17813] = 1'b0;
assign COL[17814] = 1'b0;
assign COL[17815] = 1'b0;
assign COL[17816] = 1'b0;
assign COL[17817] = 1'b0;
assign COL[17818] = 1'b0;
assign COL[17819] = 1'b0;
assign COL[17820] = 1'b0;
assign COL[17821] = 1'b0;
assign COL[17822] = 1'b0;
assign COL[17823] = 1'b0;
assign COL[17824] = 1'b0;
assign COL[17825] = 1'b0;
assign COL[17826] = 1'b0;
assign COL[17827] = 1'b0;
assign COL[17828] = 1'b0;
assign COL[17829] = 1'b0;
assign COL[17830] = 1'b0;
assign COL[17831] = 1'b0;
assign COL[17832] = 1'b0;
assign COL[17833] = 1'b0;
assign COL[17834] = 1'b0;
assign COL[17835] = 1'b0;
assign COL[17836] = 1'b0;
assign COL[17837] = 1'b0;
assign COL[17838] = 1'b0;
assign COL[17839] = 1'b0;
assign COL[17840] = 1'b0;
assign COL[17841] = 1'b0;
assign COL[17842] = 1'b0;
assign COL[17843] = 1'b0;
assign COL[17844] = 1'b0;
assign COL[17845] = 1'b0;
assign COL[17846] = 1'b0;
assign COL[17847] = 1'b0;
assign COL[17848] = 1'b0;
assign COL[17849] = 1'b0;
assign COL[17850] = 1'b0;
assign COL[17851] = 1'b0;
assign COL[17852] = 1'b0;
assign COL[17853] = 1'b0;
assign COL[17854] = 1'b0;
assign COL[17855] = 1'b0;
assign COL[17856] = 1'b0;
assign COL[17857] = 1'b0;
assign COL[17858] = 1'b0;
assign COL[17859] = 1'b0;
assign COL[17860] = 1'b0;
assign COL[17861] = 1'b0;
assign COL[17862] = 1'b0;
assign COL[17863] = 1'b0;
assign COL[17864] = 1'b0;
assign COL[17865] = 1'b0;
assign COL[17866] = 1'b0;
assign COL[17867] = 1'b0;
assign COL[17868] = 1'b0;
assign COL[17869] = 1'b0;
assign COL[17870] = 1'b0;
assign COL[17871] = 1'b0;
assign COL[17872] = 1'b0;
assign COL[17873] = 1'b0;
assign COL[17874] = 1'b0;
assign COL[17875] = 1'b0;
assign COL[17876] = 1'b0;
assign COL[17877] = 1'b0;
assign COL[17878] = 1'b0;
assign COL[17879] = 1'b0;
assign COL[17880] = 1'b0;
assign COL[17881] = 1'b0;
assign COL[17882] = 1'b0;
assign COL[17883] = 1'b0;
assign COL[17884] = 1'b0;
assign COL[17885] = 1'b0;
assign COL[17886] = 1'b0;
assign COL[17887] = 1'b0;
assign COL[17888] = 1'b0;
assign COL[17889] = 1'b0;
assign COL[17890] = 1'b0;
assign COL[17891] = 1'b0;
assign COL[17892] = 1'b0;
assign COL[17893] = 1'b0;
assign COL[17894] = 1'b0;
assign COL[17895] = 1'b0;
assign COL[17896] = 1'b0;
assign COL[17897] = 1'b0;
assign COL[17898] = 1'b0;
assign COL[17899] = 1'b0;
assign COL[17900] = 1'b0;
assign COL[17901] = 1'b0;
assign COL[17902] = 1'b0;
assign COL[17903] = 1'b0;
assign COL[17904] = 1'b0;
assign COL[17905] = 1'b0;
assign COL[17906] = 1'b0;
assign COL[17907] = 1'b0;
assign COL[17908] = 1'b0;
assign COL[17909] = 1'b0;
assign COL[17910] = 1'b0;
assign COL[17911] = 1'b0;
assign COL[17912] = 1'b0;
assign COL[17913] = 1'b0;
assign COL[17914] = 1'b0;
assign COL[17915] = 1'b0;
assign COL[17916] = 1'b0;
assign COL[17917] = 1'b0;
assign COL[17918] = 1'b0;
assign COL[17919] = 1'b0;
assign COL[17920] = 1'b0;
assign COL[17921] = 1'b0;
assign COL[17922] = 1'b0;
assign COL[17923] = 1'b0;
assign COL[17924] = 1'b0;
assign COL[17925] = 1'b0;
assign COL[17926] = 1'b0;
assign COL[17927] = 1'b0;
assign COL[17928] = 1'b0;
assign COL[17929] = 1'b0;
assign COL[17930] = 1'b0;
assign COL[17931] = 1'b0;
assign COL[17932] = 1'b0;
assign COL[17933] = 1'b0;
assign COL[17934] = 1'b0;
assign COL[17935] = 1'b0;
assign COL[17936] = 1'b0;
assign COL[17937] = 1'b0;
assign COL[17938] = 1'b0;
assign COL[17939] = 1'b0;
assign COL[17940] = 1'b0;
assign COL[17941] = 1'b0;
assign COL[17942] = 1'b0;
assign COL[17943] = 1'b0;
assign COL[17944] = 1'b0;
assign COL[17945] = 1'b0;
assign COL[17946] = 1'b0;
assign COL[17947] = 1'b0;
assign COL[17948] = 1'b0;
assign COL[17949] = 1'b0;
assign COL[17950] = 1'b0;
assign COL[17951] = 1'b0;
assign COL[17952] = 1'b0;
assign COL[17953] = 1'b0;
assign COL[17954] = 1'b0;
assign COL[17955] = 1'b0;
assign COL[17956] = 1'b0;
assign COL[17957] = 1'b0;
assign COL[17958] = 1'b0;
assign COL[17959] = 1'b0;
assign COL[17960] = 1'b0;
assign COL[17961] = 1'b0;
assign COL[17962] = 1'b0;
assign COL[17963] = 1'b0;
assign COL[17964] = 1'b0;
assign COL[17965] = 1'b0;
assign COL[17966] = 1'b0;
assign COL[17967] = 1'b0;
assign COL[17968] = 1'b0;
assign COL[17969] = 1'b0;
assign COL[17970] = 1'b0;
assign COL[17971] = 1'b0;
assign COL[17972] = 1'b0;
assign COL[17973] = 1'b0;
assign COL[17974] = 1'b0;
assign COL[17975] = 1'b0;
assign COL[17976] = 1'b0;
assign COL[17977] = 1'b0;
assign COL[17978] = 1'b0;
assign COL[17979] = 1'b0;
assign COL[17980] = 1'b0;
assign COL[17981] = 1'b0;
assign COL[17982] = 1'b0;
assign COL[17983] = 1'b0;
assign COL[17984] = 1'b0;
assign COL[17985] = 1'b0;
assign COL[17986] = 1'b0;
assign COL[17987] = 1'b0;
assign COL[17988] = 1'b0;
assign COL[17989] = 1'b0;
assign COL[17990] = 1'b0;
assign COL[17991] = 1'b0;
assign COL[17992] = 1'b0;
assign COL[17993] = 1'b0;
assign COL[17994] = 1'b0;
assign COL[17995] = 1'b0;
assign COL[17996] = 1'b0;
assign COL[17997] = 1'b0;
assign COL[17998] = 1'b0;
assign COL[17999] = 1'b0;
assign COL[18000] = 1'b0;
assign COL[18001] = 1'b0;
assign COL[18002] = 1'b0;
assign COL[18003] = 1'b0;
assign COL[18004] = 1'b0;
assign COL[18005] = 1'b0;
assign COL[18006] = 1'b0;
assign COL[18007] = 1'b0;
assign COL[18008] = 1'b0;
assign COL[18009] = 1'b0;
assign COL[18010] = 1'b0;
assign COL[18011] = 1'b0;
assign COL[18012] = 1'b0;
assign COL[18013] = 1'b0;
assign COL[18014] = 1'b0;
assign COL[18015] = 1'b0;
assign COL[18016] = 1'b0;
assign COL[18017] = 1'b0;
assign COL[18018] = 1'b0;
assign COL[18019] = 1'b0;
assign COL[18020] = 1'b0;
assign COL[18021] = 1'b0;
assign COL[18022] = 1'b0;
assign COL[18023] = 1'b0;
assign COL[18024] = 1'b0;
assign COL[18025] = 1'b0;
assign COL[18026] = 1'b0;
assign COL[18027] = 1'b0;
assign COL[18028] = 1'b0;
assign COL[18029] = 1'b0;
assign COL[18030] = 1'b0;
assign COL[18031] = 1'b0;
assign COL[18032] = 1'b0;
assign COL[18033] = 1'b0;
assign COL[18034] = 1'b0;
assign COL[18035] = 1'b0;
assign COL[18036] = 1'b0;
assign COL[18037] = 1'b0;
assign COL[18038] = 1'b0;
assign COL[18039] = 1'b0;
assign COL[18040] = 1'b0;
assign COL[18041] = 1'b0;
assign COL[18042] = 1'b0;
assign COL[18043] = 1'b0;
assign COL[18044] = 1'b0;
assign COL[18045] = 1'b0;
assign COL[18046] = 1'b0;
assign COL[18047] = 1'b0;
assign COL[18048] = 1'b0;
assign COL[18049] = 1'b0;
assign COL[18050] = 1'b0;
assign COL[18051] = 1'b0;
assign COL[18052] = 1'b0;
assign COL[18053] = 1'b0;
assign COL[18054] = 1'b0;
assign COL[18055] = 1'b0;
assign COL[18056] = 1'b0;
assign COL[18057] = 1'b0;
assign COL[18058] = 1'b0;
assign COL[18059] = 1'b0;
assign COL[18060] = 1'b0;
assign COL[18061] = 1'b0;
assign COL[18062] = 1'b0;
assign COL[18063] = 1'b0;
assign COL[18064] = 1'b0;
assign COL[18065] = 1'b0;
assign COL[18066] = 1'b0;
assign COL[18067] = 1'b0;
assign COL[18068] = 1'b0;
assign COL[18069] = 1'b0;
assign COL[18070] = 1'b0;
assign COL[18071] = 1'b0;
assign COL[18072] = 1'b0;
assign COL[18073] = 1'b0;
assign COL[18074] = 1'b0;
assign COL[18075] = 1'b0;
assign COL[18076] = 1'b0;
assign COL[18077] = 1'b0;
assign COL[18078] = 1'b0;
assign COL[18079] = 1'b0;
assign COL[18080] = 1'b0;
assign COL[18081] = 1'b0;
assign COL[18082] = 1'b0;
assign COL[18083] = 1'b0;
assign COL[18084] = 1'b0;
assign COL[18085] = 1'b0;
assign COL[18086] = 1'b0;
assign COL[18087] = 1'b0;
assign COL[18088] = 1'b0;
assign COL[18089] = 1'b0;
assign COL[18090] = 1'b0;
assign COL[18091] = 1'b0;
assign COL[18092] = 1'b0;
assign COL[18093] = 1'b0;
assign COL[18094] = 1'b0;
assign COL[18095] = 1'b0;
assign COL[18096] = 1'b0;
assign COL[18097] = 1'b0;
assign COL[18098] = 1'b0;
assign COL[18099] = 1'b0;
assign COL[18100] = 1'b0;
assign COL[18101] = 1'b0;
assign COL[18102] = 1'b0;
assign COL[18103] = 1'b0;
assign COL[18104] = 1'b0;
assign COL[18105] = 1'b0;
assign COL[18106] = 1'b0;
assign COL[18107] = 1'b0;
assign COL[18108] = 1'b0;
assign COL[18109] = 1'b0;
assign COL[18110] = 1'b0;
assign COL[18111] = 1'b0;
assign COL[18112] = 1'b0;
assign COL[18113] = 1'b0;
assign COL[18114] = 1'b0;
assign COL[18115] = 1'b0;
assign COL[18116] = 1'b0;
assign COL[18117] = 1'b0;
assign COL[18118] = 1'b0;
assign COL[18119] = 1'b0;
assign COL[18120] = 1'b0;
assign COL[18121] = 1'b0;
assign COL[18122] = 1'b0;
assign COL[18123] = 1'b0;
assign COL[18124] = 1'b0;
assign COL[18125] = 1'b0;
assign COL[18126] = 1'b0;
assign COL[18127] = 1'b0;
assign COL[18128] = 1'b0;
assign COL[18129] = 1'b0;
assign COL[18130] = 1'b0;
assign COL[18131] = 1'b0;
assign COL[18132] = 1'b0;
assign COL[18133] = 1'b0;
assign COL[18134] = 1'b0;
assign COL[18135] = 1'b0;
assign COL[18136] = 1'b0;
assign COL[18137] = 1'b0;
assign COL[18138] = 1'b0;
assign COL[18139] = 1'b0;
assign COL[18140] = 1'b0;
assign COL[18141] = 1'b0;
assign COL[18142] = 1'b0;
assign COL[18143] = 1'b0;
assign COL[18144] = 1'b0;
assign COL[18145] = 1'b0;
assign COL[18146] = 1'b0;
assign COL[18147] = 1'b0;
assign COL[18148] = 1'b0;
assign COL[18149] = 1'b0;
assign COL[18150] = 1'b0;
assign COL[18151] = 1'b0;
assign COL[18152] = 1'b0;
assign COL[18153] = 1'b0;
assign COL[18154] = 1'b0;
assign COL[18155] = 1'b0;
assign COL[18156] = 1'b0;
assign COL[18157] = 1'b0;
assign COL[18158] = 1'b0;
assign COL[18159] = 1'b0;
assign COL[18160] = 1'b0;
assign COL[18161] = 1'b0;
assign COL[18162] = 1'b0;
assign COL[18163] = 1'b0;
assign COL[18164] = 1'b0;
assign COL[18165] = 1'b0;
assign COL[18166] = 1'b0;
assign COL[18167] = 1'b0;
assign COL[18168] = 1'b0;
assign COL[18169] = 1'b0;
assign COL[18170] = 1'b0;
assign COL[18171] = 1'b0;
assign COL[18172] = 1'b0;
assign COL[18173] = 1'b0;
assign COL[18174] = 1'b0;
assign COL[18175] = 1'b0;
assign COL[18176] = 1'b0;
assign COL[18177] = 1'b0;
assign COL[18178] = 1'b0;
assign COL[18179] = 1'b0;
assign COL[18180] = 1'b0;
assign COL[18181] = 1'b0;
assign COL[18182] = 1'b0;
assign COL[18183] = 1'b0;
assign COL[18184] = 1'b0;
assign COL[18185] = 1'b0;
assign COL[18186] = 1'b0;
assign COL[18187] = 1'b0;
assign COL[18188] = 1'b0;
assign COL[18189] = 1'b0;
assign COL[18190] = 1'b0;
assign COL[18191] = 1'b0;
assign COL[18192] = 1'b0;
assign COL[18193] = 1'b0;
assign COL[18194] = 1'b0;
assign COL[18195] = 1'b0;
assign COL[18196] = 1'b0;
assign COL[18197] = 1'b0;
assign COL[18198] = 1'b0;
assign COL[18199] = 1'b0;
assign COL[18200] = 1'b0;
assign COL[18201] = 1'b0;
assign COL[18202] = 1'b0;
assign COL[18203] = 1'b0;
assign COL[18204] = 1'b0;
assign COL[18205] = 1'b0;
assign COL[18206] = 1'b0;
assign COL[18207] = 1'b0;
assign COL[18208] = 1'b0;
assign COL[18209] = 1'b0;
assign COL[18210] = 1'b0;
assign COL[18211] = 1'b0;
assign COL[18212] = 1'b0;
assign COL[18213] = 1'b0;
assign COL[18214] = 1'b0;
assign COL[18215] = 1'b0;
assign COL[18216] = 1'b0;
assign COL[18217] = 1'b0;
assign COL[18218] = 1'b0;
assign COL[18219] = 1'b0;
assign COL[18220] = 1'b0;
assign COL[18221] = 1'b0;
assign COL[18222] = 1'b0;
assign COL[18223] = 1'b0;
assign COL[18224] = 1'b0;
assign COL[18225] = 1'b0;
assign COL[18226] = 1'b0;
assign COL[18227] = 1'b0;
assign COL[18228] = 1'b0;
assign COL[18229] = 1'b0;
assign COL[18230] = 1'b0;
assign COL[18231] = 1'b0;
assign COL[18232] = 1'b0;
assign COL[18233] = 1'b0;
assign COL[18234] = 1'b0;
assign COL[18235] = 1'b0;
assign COL[18236] = 1'b0;
assign COL[18237] = 1'b0;
assign COL[18238] = 1'b0;
assign COL[18239] = 1'b0;
assign COL[18240] = 1'b0;
assign COL[18241] = 1'b0;
assign COL[18242] = 1'b0;
assign COL[18243] = 1'b0;
assign COL[18244] = 1'b0;
assign COL[18245] = 1'b0;
assign COL[18246] = 1'b0;
assign COL[18247] = 1'b0;
assign COL[18248] = 1'b0;
assign COL[18249] = 1'b0;
assign COL[18250] = 1'b0;
assign COL[18251] = 1'b0;
assign COL[18252] = 1'b0;
assign COL[18253] = 1'b0;
assign COL[18254] = 1'b0;
assign COL[18255] = 1'b0;
assign COL[18256] = 1'b0;
assign COL[18257] = 1'b0;
assign COL[18258] = 1'b0;
assign COL[18259] = 1'b0;
assign COL[18260] = 1'b0;
assign COL[18261] = 1'b0;
assign COL[18262] = 1'b0;
assign COL[18263] = 1'b0;
assign COL[18264] = 1'b0;
assign COL[18265] = 1'b0;
assign COL[18266] = 1'b0;
assign COL[18267] = 1'b0;
assign COL[18268] = 1'b0;
assign COL[18269] = 1'b0;
assign COL[18270] = 1'b0;
assign COL[18271] = 1'b0;
assign COL[18272] = 1'b0;
assign COL[18273] = 1'b0;
assign COL[18274] = 1'b0;
assign COL[18275] = 1'b0;
assign COL[18276] = 1'b0;
assign COL[18277] = 1'b0;
assign COL[18278] = 1'b0;
assign COL[18279] = 1'b0;
assign COL[18280] = 1'b0;
assign COL[18281] = 1'b0;
assign COL[18282] = 1'b0;
assign COL[18283] = 1'b0;
assign COL[18284] = 1'b0;
assign COL[18285] = 1'b0;
assign COL[18286] = 1'b0;
assign COL[18287] = 1'b0;
assign COL[18288] = 1'b0;
assign COL[18289] = 1'b0;
assign COL[18290] = 1'b0;
assign COL[18291] = 1'b0;
assign COL[18292] = 1'b0;
assign COL[18293] = 1'b0;
assign COL[18294] = 1'b0;
assign COL[18295] = 1'b0;
assign COL[18296] = 1'b0;
assign COL[18297] = 1'b0;
assign COL[18298] = 1'b0;
assign COL[18299] = 1'b0;
assign COL[18300] = 1'b0;
assign COL[18301] = 1'b0;
assign COL[18302] = 1'b0;
assign COL[18303] = 1'b0;
assign COL[18304] = 1'b0;
assign COL[18305] = 1'b0;
assign COL[18306] = 1'b0;
assign COL[18307] = 1'b0;
assign COL[18308] = 1'b0;
assign COL[18309] = 1'b0;
assign COL[18310] = 1'b0;
assign COL[18311] = 1'b0;
assign COL[18312] = 1'b0;
assign COL[18313] = 1'b0;
assign COL[18314] = 1'b0;
assign COL[18315] = 1'b0;
assign COL[18316] = 1'b0;
assign COL[18317] = 1'b0;
assign COL[18318] = 1'b0;
assign COL[18319] = 1'b0;
assign COL[18320] = 1'b0;
assign COL[18321] = 1'b0;
assign COL[18322] = 1'b0;
assign COL[18323] = 1'b0;
assign COL[18324] = 1'b0;
assign COL[18325] = 1'b0;
assign COL[18326] = 1'b0;
assign COL[18327] = 1'b0;
assign COL[18328] = 1'b0;
assign COL[18329] = 1'b0;
assign COL[18330] = 1'b0;
assign COL[18331] = 1'b0;
assign COL[18332] = 1'b0;
assign COL[18333] = 1'b0;
assign COL[18334] = 1'b0;
assign COL[18335] = 1'b0;
assign COL[18336] = 1'b0;
assign COL[18337] = 1'b0;
assign COL[18338] = 1'b0;
assign COL[18339] = 1'b0;
assign COL[18340] = 1'b0;
assign COL[18341] = 1'b0;
assign COL[18342] = 1'b0;
assign COL[18343] = 1'b0;
assign COL[18344] = 1'b0;
assign COL[18345] = 1'b0;
assign COL[18346] = 1'b0;
assign COL[18347] = 1'b0;
assign COL[18348] = 1'b0;
assign COL[18349] = 1'b0;
assign COL[18350] = 1'b0;
assign COL[18351] = 1'b0;
assign COL[18352] = 1'b0;
assign COL[18353] = 1'b0;
assign COL[18354] = 1'b0;
assign COL[18355] = 1'b0;
assign COL[18356] = 1'b0;
assign COL[18357] = 1'b0;
assign COL[18358] = 1'b0;
assign COL[18359] = 1'b0;
assign COL[18360] = 1'b0;
assign COL[18361] = 1'b0;
assign COL[18362] = 1'b0;
assign COL[18363] = 1'b0;
assign COL[18364] = 1'b0;
assign COL[18365] = 1'b0;
assign COL[18366] = 1'b0;
assign COL[18367] = 1'b0;
assign COL[18368] = 1'b0;
assign COL[18369] = 1'b0;
assign COL[18370] = 1'b0;
assign COL[18371] = 1'b0;
assign COL[18372] = 1'b0;
assign COL[18373] = 1'b0;
assign COL[18374] = 1'b0;
assign COL[18375] = 1'b0;
assign COL[18376] = 1'b0;
assign COL[18377] = 1'b0;
assign COL[18378] = 1'b0;
assign COL[18379] = 1'b0;
assign COL[18380] = 1'b0;
assign COL[18381] = 1'b0;
assign COL[18382] = 1'b0;
assign COL[18383] = 1'b0;
assign COL[18384] = 1'b0;
assign COL[18385] = 1'b0;
assign COL[18386] = 1'b0;
assign COL[18387] = 1'b0;
assign COL[18388] = 1'b0;
assign COL[18389] = 1'b0;
assign COL[18390] = 1'b0;
assign COL[18391] = 1'b0;
assign COL[18392] = 1'b0;
assign COL[18393] = 1'b0;
assign COL[18394] = 1'b0;
assign COL[18395] = 1'b0;
assign COL[18396] = 1'b0;
assign COL[18397] = 1'b0;
assign COL[18398] = 1'b0;
assign COL[18399] = 1'b0;
assign COL[18400] = 1'b0;
assign COL[18401] = 1'b0;
assign COL[18402] = 1'b0;
assign COL[18403] = 1'b0;
assign COL[18404] = 1'b0;
assign COL[18405] = 1'b0;
assign COL[18406] = 1'b0;
assign COL[18407] = 1'b0;
assign COL[18408] = 1'b0;
assign COL[18409] = 1'b0;
assign COL[18410] = 1'b0;
assign COL[18411] = 1'b0;
assign COL[18412] = 1'b0;
assign COL[18413] = 1'b0;
assign COL[18414] = 1'b0;
assign COL[18415] = 1'b0;
assign COL[18416] = 1'b0;
assign COL[18417] = 1'b0;
assign COL[18418] = 1'b0;
assign COL[18419] = 1'b0;
assign COL[18420] = 1'b0;
assign COL[18421] = 1'b0;
assign COL[18422] = 1'b0;
assign COL[18423] = 1'b0;
assign COL[18424] = 1'b0;
assign COL[18425] = 1'b0;
assign COL[18426] = 1'b0;
assign COL[18427] = 1'b0;
assign COL[18428] = 1'b0;
assign COL[18429] = 1'b0;
assign COL[18430] = 1'b0;
assign COL[18431] = 1'b0;
assign COL[18432] = 1'b0;
assign COL[18433] = 1'b0;
assign COL[18434] = 1'b0;
assign COL[18435] = 1'b0;
assign COL[18436] = 1'b0;
assign COL[18437] = 1'b0;
assign COL[18438] = 1'b0;
assign COL[18439] = 1'b0;
assign COL[18440] = 1'b0;
assign COL[18441] = 1'b0;
assign COL[18442] = 1'b0;
assign COL[18443] = 1'b0;
assign COL[18444] = 1'b0;
assign COL[18445] = 1'b0;
assign COL[18446] = 1'b0;
assign COL[18447] = 1'b0;
assign COL[18448] = 1'b0;
assign COL[18449] = 1'b0;
assign COL[18450] = 1'b0;
assign COL[18451] = 1'b0;
assign COL[18452] = 1'b0;
assign COL[18453] = 1'b0;
assign COL[18454] = 1'b0;
assign COL[18455] = 1'b0;
assign COL[18456] = 1'b0;
assign COL[18457] = 1'b0;
assign COL[18458] = 1'b0;
assign COL[18459] = 1'b0;
assign COL[18460] = 1'b0;
assign COL[18461] = 1'b0;
assign COL[18462] = 1'b0;
assign COL[18463] = 1'b0;
assign COL[18464] = 1'b0;
assign COL[18465] = 1'b0;
assign COL[18466] = 1'b0;
assign COL[18467] = 1'b0;
assign COL[18468] = 1'b0;
assign COL[18469] = 1'b0;
assign COL[18470] = 1'b0;
assign COL[18471] = 1'b0;
assign COL[18472] = 1'b0;
assign COL[18473] = 1'b0;
assign COL[18474] = 1'b0;
assign COL[18475] = 1'b0;
assign COL[18476] = 1'b0;
assign COL[18477] = 1'b0;
assign COL[18478] = 1'b0;
assign COL[18479] = 1'b0;
assign COL[18480] = 1'b0;
assign COL[18481] = 1'b0;
assign COL[18482] = 1'b0;
assign COL[18483] = 1'b0;
assign COL[18484] = 1'b0;
assign COL[18485] = 1'b0;
assign COL[18486] = 1'b0;
assign COL[18487] = 1'b0;
assign COL[18488] = 1'b0;
assign COL[18489] = 1'b0;
assign COL[18490] = 1'b0;
assign COL[18491] = 1'b0;
assign COL[18492] = 1'b0;
assign COL[18493] = 1'b0;
assign COL[18494] = 1'b0;
assign COL[18495] = 1'b0;
assign COL[18496] = 1'b0;
assign COL[18497] = 1'b0;
assign COL[18498] = 1'b0;
assign COL[18499] = 1'b0;
assign COL[18500] = 1'b0;
assign COL[18501] = 1'b0;
assign COL[18502] = 1'b0;
assign COL[18503] = 1'b0;
assign COL[18504] = 1'b0;
assign COL[18505] = 1'b0;
assign COL[18506] = 1'b0;
assign COL[18507] = 1'b0;
assign COL[18508] = 1'b0;
assign COL[18509] = 1'b0;
assign COL[18510] = 1'b0;
assign COL[18511] = 1'b0;
assign COL[18512] = 1'b0;
assign COL[18513] = 1'b0;
assign COL[18514] = 1'b0;
assign COL[18515] = 1'b0;
assign COL[18516] = 1'b0;
assign COL[18517] = 1'b0;
assign COL[18518] = 1'b0;
assign COL[18519] = 1'b0;
assign COL[18520] = 1'b0;
assign COL[18521] = 1'b0;
assign COL[18522] = 1'b0;
assign COL[18523] = 1'b0;
assign COL[18524] = 1'b0;
assign COL[18525] = 1'b0;
assign COL[18526] = 1'b0;
assign COL[18527] = 1'b0;
assign COL[18528] = 1'b0;
assign COL[18529] = 1'b0;
assign COL[18530] = 1'b0;
assign COL[18531] = 1'b0;
assign COL[18532] = 1'b0;
assign COL[18533] = 1'b0;
assign COL[18534] = 1'b0;
assign COL[18535] = 1'b0;
assign COL[18536] = 1'b0;
assign COL[18537] = 1'b0;
assign COL[18538] = 1'b0;
assign COL[18539] = 1'b0;
assign COL[18540] = 1'b0;
assign COL[18541] = 1'b0;
assign COL[18542] = 1'b0;
assign COL[18543] = 1'b0;
assign COL[18544] = 1'b0;
assign COL[18545] = 1'b0;
assign COL[18546] = 1'b0;
assign COL[18547] = 1'b0;
assign COL[18548] = 1'b0;
assign COL[18549] = 1'b0;
assign COL[18550] = 1'b0;
assign COL[18551] = 1'b0;
assign COL[18552] = 1'b0;
assign COL[18553] = 1'b0;
assign COL[18554] = 1'b0;
assign COL[18555] = 1'b0;
assign COL[18556] = 1'b0;
assign COL[18557] = 1'b0;
assign COL[18558] = 1'b0;
assign COL[18559] = 1'b0;
assign COL[18560] = 1'b0;
assign COL[18561] = 1'b0;
assign COL[18562] = 1'b0;
assign COL[18563] = 1'b0;
assign COL[18564] = 1'b0;
assign COL[18565] = 1'b0;
assign COL[18566] = 1'b0;
assign COL[18567] = 1'b0;
assign COL[18568] = 1'b0;
assign COL[18569] = 1'b0;
assign COL[18570] = 1'b0;
assign COL[18571] = 1'b0;
assign COL[18572] = 1'b0;
assign COL[18573] = 1'b0;
assign COL[18574] = 1'b0;
assign COL[18575] = 1'b0;
assign COL[18576] = 1'b0;
assign COL[18577] = 1'b0;
assign COL[18578] = 1'b0;
assign COL[18579] = 1'b0;
assign COL[18580] = 1'b0;
assign COL[18581] = 1'b0;
assign COL[18582] = 1'b0;
assign COL[18583] = 1'b0;
assign COL[18584] = 1'b0;
assign COL[18585] = 1'b0;
assign COL[18586] = 1'b0;
assign COL[18587] = 1'b0;
assign COL[18588] = 1'b0;
assign COL[18589] = 1'b0;
assign COL[18590] = 1'b0;
assign COL[18591] = 1'b0;
assign COL[18592] = 1'b0;
assign COL[18593] = 1'b0;
assign COL[18594] = 1'b0;
assign COL[18595] = 1'b0;
assign COL[18596] = 1'b0;
assign COL[18597] = 1'b0;
assign COL[18598] = 1'b0;
assign COL[18599] = 1'b0;
assign COL[18600] = 1'b0;
assign COL[18601] = 1'b0;
assign COL[18602] = 1'b0;
assign COL[18603] = 1'b0;
assign COL[18604] = 1'b0;
assign COL[18605] = 1'b0;
assign COL[18606] = 1'b0;
assign COL[18607] = 1'b0;
assign COL[18608] = 1'b0;
assign COL[18609] = 1'b0;
assign COL[18610] = 1'b0;
assign COL[18611] = 1'b0;
assign COL[18612] = 1'b0;
assign COL[18613] = 1'b0;
assign COL[18614] = 1'b0;
assign COL[18615] = 1'b0;
assign COL[18616] = 1'b0;
assign COL[18617] = 1'b0;
assign COL[18618] = 1'b0;
assign COL[18619] = 1'b0;
assign COL[18620] = 1'b0;
assign COL[18621] = 1'b0;
assign COL[18622] = 1'b0;
assign COL[18623] = 1'b0;
assign COL[18624] = 1'b0;
assign COL[18625] = 1'b0;
assign COL[18626] = 1'b0;
assign COL[18627] = 1'b0;
assign COL[18628] = 1'b0;
assign COL[18629] = 1'b0;
assign COL[18630] = 1'b0;
assign COL[18631] = 1'b0;
assign COL[18632] = 1'b0;
assign COL[18633] = 1'b0;
assign COL[18634] = 1'b0;
assign COL[18635] = 1'b0;
assign COL[18636] = 1'b0;
assign COL[18637] = 1'b0;
assign COL[18638] = 1'b0;
assign COL[18639] = 1'b0;
assign COL[18640] = 1'b0;
assign COL[18641] = 1'b0;
assign COL[18642] = 1'b0;
assign COL[18643] = 1'b0;
assign COL[18644] = 1'b0;
assign COL[18645] = 1'b0;
assign COL[18646] = 1'b0;
assign COL[18647] = 1'b0;
assign COL[18648] = 1'b0;
assign COL[18649] = 1'b0;
assign COL[18650] = 1'b0;
assign COL[18651] = 1'b0;
assign COL[18652] = 1'b0;
assign COL[18653] = 1'b0;
assign COL[18654] = 1'b0;
assign COL[18655] = 1'b0;
assign COL[18656] = 1'b0;
assign COL[18657] = 1'b0;
assign COL[18658] = 1'b0;
assign COL[18659] = 1'b0;
assign COL[18660] = 1'b0;
assign COL[18661] = 1'b0;
assign COL[18662] = 1'b0;
assign COL[18663] = 1'b0;
assign COL[18664] = 1'b0;
assign COL[18665] = 1'b0;
assign COL[18666] = 1'b0;
assign COL[18667] = 1'b0;
assign COL[18668] = 1'b0;
assign COL[18669] = 1'b0;
assign COL[18670] = 1'b0;
assign COL[18671] = 1'b0;
assign COL[18672] = 1'b0;
assign COL[18673] = 1'b0;
assign COL[18674] = 1'b0;
assign COL[18675] = 1'b0;
assign COL[18676] = 1'b0;
assign COL[18677] = 1'b0;
assign COL[18678] = 1'b0;
assign COL[18679] = 1'b0;
assign COL[18680] = 1'b0;
assign COL[18681] = 1'b0;
assign COL[18682] = 1'b0;
assign COL[18683] = 1'b0;
assign COL[18684] = 1'b0;
assign COL[18685] = 1'b0;
assign COL[18686] = 1'b0;
assign COL[18687] = 1'b0;
assign COL[18688] = 1'b0;
assign COL[18689] = 1'b0;
assign COL[18690] = 1'b0;
assign COL[18691] = 1'b0;
assign COL[18692] = 1'b0;
assign COL[18693] = 1'b0;
assign COL[18694] = 1'b0;
assign COL[18695] = 1'b0;
assign COL[18696] = 1'b0;
assign COL[18697] = 1'b0;
assign COL[18698] = 1'b0;
assign COL[18699] = 1'b0;
assign COL[18700] = 1'b0;
assign COL[18701] = 1'b0;
assign COL[18702] = 1'b0;
assign COL[18703] = 1'b0;
assign COL[18704] = 1'b0;
assign COL[18705] = 1'b0;
assign COL[18706] = 1'b0;
assign COL[18707] = 1'b0;
assign COL[18708] = 1'b0;
assign COL[18709] = 1'b0;
assign COL[18710] = 1'b0;
assign COL[18711] = 1'b0;
assign COL[18712] = 1'b0;
assign COL[18713] = 1'b0;
assign COL[18714] = 1'b0;
assign COL[18715] = 1'b0;
assign COL[18716] = 1'b0;
assign COL[18717] = 1'b0;
assign COL[18718] = 1'b0;
assign COL[18719] = 1'b0;
assign COL[18720] = 1'b0;
assign COL[18721] = 1'b0;
assign COL[18722] = 1'b0;
assign COL[18723] = 1'b0;
assign COL[18724] = 1'b0;
assign COL[18725] = 1'b0;
assign COL[18726] = 1'b0;
assign COL[18727] = 1'b0;
assign COL[18728] = 1'b0;
assign COL[18729] = 1'b0;
assign COL[18730] = 1'b0;
assign COL[18731] = 1'b0;
assign COL[18732] = 1'b0;
assign COL[18733] = 1'b0;
assign COL[18734] = 1'b0;
assign COL[18735] = 1'b0;
assign COL[18736] = 1'b0;
assign COL[18737] = 1'b0;
assign COL[18738] = 1'b0;
assign COL[18739] = 1'b0;
assign COL[18740] = 1'b0;
assign COL[18741] = 1'b0;
assign COL[18742] = 1'b0;
assign COL[18743] = 1'b0;
assign COL[18744] = 1'b0;
assign COL[18745] = 1'b0;
assign COL[18746] = 1'b0;
assign COL[18747] = 1'b0;
assign COL[18748] = 1'b0;
assign COL[18749] = 1'b0;
assign COL[18750] = 1'b0;
assign COL[18751] = 1'b0;
assign COL[18752] = 1'b0;
assign COL[18753] = 1'b0;
assign COL[18754] = 1'b0;
assign COL[18755] = 1'b0;
assign COL[18756] = 1'b0;
assign COL[18757] = 1'b0;
assign COL[18758] = 1'b0;
assign COL[18759] = 1'b0;
assign COL[18760] = 1'b0;
assign COL[18761] = 1'b0;
assign COL[18762] = 1'b0;
assign COL[18763] = 1'b0;
assign COL[18764] = 1'b0;
assign COL[18765] = 1'b0;
assign COL[18766] = 1'b0;
assign COL[18767] = 1'b0;
assign COL[18768] = 1'b0;
assign COL[18769] = 1'b0;
assign COL[18770] = 1'b0;
assign COL[18771] = 1'b0;
assign COL[18772] = 1'b0;
assign COL[18773] = 1'b0;
assign COL[18774] = 1'b0;
assign COL[18775] = 1'b0;
assign COL[18776] = 1'b0;
assign COL[18777] = 1'b0;
assign COL[18778] = 1'b0;
assign COL[18779] = 1'b0;
assign COL[18780] = 1'b0;
assign COL[18781] = 1'b0;
assign COL[18782] = 1'b0;
assign COL[18783] = 1'b0;
assign COL[18784] = 1'b0;
assign COL[18785] = 1'b0;
assign COL[18786] = 1'b0;
assign COL[18787] = 1'b0;
assign COL[18788] = 1'b0;
assign COL[18789] = 1'b0;
assign COL[18790] = 1'b0;
assign COL[18791] = 1'b0;
assign COL[18792] = 1'b0;
assign COL[18793] = 1'b0;
assign COL[18794] = 1'b0;
assign COL[18795] = 1'b0;
assign COL[18796] = 1'b0;
assign COL[18797] = 1'b0;
assign COL[18798] = 1'b0;
assign COL[18799] = 1'b0;
assign COL[18800] = 1'b0;
assign COL[18801] = 1'b0;
assign COL[18802] = 1'b0;
assign COL[18803] = 1'b0;
assign COL[18804] = 1'b0;
assign COL[18805] = 1'b0;
assign COL[18806] = 1'b0;
assign COL[18807] = 1'b0;
assign COL[18808] = 1'b0;
assign COL[18809] = 1'b0;
assign COL[18810] = 1'b0;
assign COL[18811] = 1'b0;
assign COL[18812] = 1'b0;
assign COL[18813] = 1'b0;
assign COL[18814] = 1'b0;
assign COL[18815] = 1'b0;
assign COL[18816] = 1'b0;
assign COL[18817] = 1'b0;
assign COL[18818] = 1'b0;
assign COL[18819] = 1'b0;
assign COL[18820] = 1'b0;
assign COL[18821] = 1'b0;
assign COL[18822] = 1'b0;
assign COL[18823] = 1'b0;
assign COL[18824] = 1'b0;
assign COL[18825] = 1'b0;
assign COL[18826] = 1'b0;
assign COL[18827] = 1'b0;
assign COL[18828] = 1'b0;
assign COL[18829] = 1'b0;
assign COL[18830] = 1'b0;
assign COL[18831] = 1'b0;
assign COL[18832] = 1'b0;
assign COL[18833] = 1'b0;
assign COL[18834] = 1'b0;
assign COL[18835] = 1'b0;
assign COL[18836] = 1'b0;
assign COL[18837] = 1'b0;
assign COL[18838] = 1'b0;
assign COL[18839] = 1'b0;
assign COL[18840] = 1'b0;
assign COL[18841] = 1'b0;
assign COL[18842] = 1'b0;
assign COL[18843] = 1'b0;
assign COL[18844] = 1'b0;
assign COL[18845] = 1'b0;
assign COL[18846] = 1'b0;
assign COL[18847] = 1'b0;
assign COL[18848] = 1'b0;
assign COL[18849] = 1'b0;
assign COL[18850] = 1'b0;
assign COL[18851] = 1'b0;
assign COL[18852] = 1'b0;
assign COL[18853] = 1'b0;
assign COL[18854] = 1'b0;
assign COL[18855] = 1'b0;
assign COL[18856] = 1'b0;
assign COL[18857] = 1'b0;
assign COL[18858] = 1'b0;
assign COL[18859] = 1'b0;
assign COL[18860] = 1'b0;
assign COL[18861] = 1'b0;
assign COL[18862] = 1'b0;
assign COL[18863] = 1'b0;
assign COL[18864] = 1'b0;
assign COL[18865] = 1'b0;
assign COL[18866] = 1'b0;
assign COL[18867] = 1'b0;
assign COL[18868] = 1'b0;
assign COL[18869] = 1'b0;
assign COL[18870] = 1'b0;
assign COL[18871] = 1'b0;
assign COL[18872] = 1'b0;
assign COL[18873] = 1'b0;
assign COL[18874] = 1'b0;
assign COL[18875] = 1'b0;
assign COL[18876] = 1'b0;
assign COL[18877] = 1'b0;
assign COL[18878] = 1'b0;
assign COL[18879] = 1'b0;
assign COL[18880] = 1'b0;
assign COL[18881] = 1'b0;
assign COL[18882] = 1'b0;
assign COL[18883] = 1'b0;
assign COL[18884] = 1'b0;
assign COL[18885] = 1'b0;
assign COL[18886] = 1'b0;
assign COL[18887] = 1'b0;
assign COL[18888] = 1'b0;
assign COL[18889] = 1'b0;
assign COL[18890] = 1'b0;
assign COL[18891] = 1'b0;
assign COL[18892] = 1'b0;
assign COL[18893] = 1'b0;
assign COL[18894] = 1'b0;
assign COL[18895] = 1'b0;
assign COL[18896] = 1'b0;
assign COL[18897] = 1'b0;
assign COL[18898] = 1'b0;
assign COL[18899] = 1'b0;
assign COL[18900] = 1'b0;
assign COL[18901] = 1'b0;
assign COL[18902] = 1'b0;
assign COL[18903] = 1'b0;
assign COL[18904] = 1'b0;
assign COL[18905] = 1'b0;
assign COL[18906] = 1'b0;
assign COL[18907] = 1'b0;
assign COL[18908] = 1'b0;
assign COL[18909] = 1'b0;
assign COL[18910] = 1'b0;
assign COL[18911] = 1'b0;
assign COL[18912] = 1'b0;
assign COL[18913] = 1'b0;
assign COL[18914] = 1'b0;
assign COL[18915] = 1'b0;
assign COL[18916] = 1'b0;
assign COL[18917] = 1'b0;
assign COL[18918] = 1'b0;
assign COL[18919] = 1'b0;
assign COL[18920] = 1'b0;
assign COL[18921] = 1'b0;
assign COL[18922] = 1'b0;
assign COL[18923] = 1'b0;
assign COL[18924] = 1'b0;
assign COL[18925] = 1'b0;
assign COL[18926] = 1'b0;
assign COL[18927] = 1'b0;
assign COL[18928] = 1'b0;
assign COL[18929] = 1'b0;
assign COL[18930] = 1'b0;
assign COL[18931] = 1'b0;
assign COL[18932] = 1'b0;
assign COL[18933] = 1'b0;
assign COL[18934] = 1'b0;
assign COL[18935] = 1'b0;
assign COL[18936] = 1'b0;
assign COL[18937] = 1'b0;
assign COL[18938] = 1'b0;
assign COL[18939] = 1'b0;
assign COL[18940] = 1'b0;
assign COL[18941] = 1'b0;
assign COL[18942] = 1'b0;
assign COL[18943] = 1'b0;
assign COL[18944] = 1'b0;
assign COL[18945] = 1'b0;
assign COL[18946] = 1'b0;
assign COL[18947] = 1'b0;
assign COL[18948] = 1'b0;
assign COL[18949] = 1'b0;
assign COL[18950] = 1'b0;
assign COL[18951] = 1'b0;
assign COL[18952] = 1'b0;
assign COL[18953] = 1'b0;
assign COL[18954] = 1'b0;
assign COL[18955] = 1'b0;
assign COL[18956] = 1'b0;
assign COL[18957] = 1'b0;
assign COL[18958] = 1'b0;
assign COL[18959] = 1'b0;
assign COL[18960] = 1'b0;
assign COL[18961] = 1'b0;
assign COL[18962] = 1'b0;
assign COL[18963] = 1'b0;
assign COL[18964] = 1'b0;
assign COL[18965] = 1'b0;
assign COL[18966] = 1'b0;
assign COL[18967] = 1'b0;
assign COL[18968] = 1'b0;
assign COL[18969] = 1'b0;
assign COL[18970] = 1'b0;
assign COL[18971] = 1'b0;
assign COL[18972] = 1'b0;
assign COL[18973] = 1'b0;
assign COL[18974] = 1'b0;
assign COL[18975] = 1'b0;
assign COL[18976] = 1'b0;
assign COL[18977] = 1'b0;
assign COL[18978] = 1'b0;
assign COL[18979] = 1'b0;
assign COL[18980] = 1'b0;
assign COL[18981] = 1'b0;
assign COL[18982] = 1'b0;
assign COL[18983] = 1'b0;
assign COL[18984] = 1'b0;
assign COL[18985] = 1'b0;
assign COL[18986] = 1'b0;
assign COL[18987] = 1'b0;
assign COL[18988] = 1'b0;
assign COL[18989] = 1'b0;
assign COL[18990] = 1'b0;
assign COL[18991] = 1'b0;
assign COL[18992] = 1'b0;
assign COL[18993] = 1'b0;
assign COL[18994] = 1'b0;
assign COL[18995] = 1'b0;
assign COL[18996] = 1'b0;
assign COL[18997] = 1'b0;
assign COL[18998] = 1'b0;
assign COL[18999] = 1'b0;
assign COL[19000] = 1'b0;
assign COL[19001] = 1'b0;
assign COL[19002] = 1'b0;
assign COL[19003] = 1'b0;
assign COL[19004] = 1'b0;
assign COL[19005] = 1'b0;
assign COL[19006] = 1'b0;
assign COL[19007] = 1'b0;
assign COL[19008] = 1'b0;
assign COL[19009] = 1'b0;
assign COL[19010] = 1'b0;
assign COL[19011] = 1'b0;
assign COL[19012] = 1'b0;
assign COL[19013] = 1'b0;
assign COL[19014] = 1'b0;
assign COL[19015] = 1'b0;
assign COL[19016] = 1'b0;
assign COL[19017] = 1'b0;
assign COL[19018] = 1'b0;
assign COL[19019] = 1'b0;
assign COL[19020] = 1'b0;
assign COL[19021] = 1'b0;
assign COL[19022] = 1'b0;
assign COL[19023] = 1'b0;
assign COL[19024] = 1'b0;
assign COL[19025] = 1'b0;
assign COL[19026] = 1'b0;
assign COL[19027] = 1'b0;
assign COL[19028] = 1'b0;
assign COL[19029] = 1'b0;
assign COL[19030] = 1'b0;
assign COL[19031] = 1'b0;
assign COL[19032] = 1'b0;
assign COL[19033] = 1'b0;
assign COL[19034] = 1'b0;
assign COL[19035] = 1'b0;
assign COL[19036] = 1'b0;
assign COL[19037] = 1'b0;
assign COL[19038] = 1'b0;
assign COL[19039] = 1'b0;
assign COL[19040] = 1'b0;
assign COL[19041] = 1'b0;
assign COL[19042] = 1'b0;
assign COL[19043] = 1'b0;
assign COL[19044] = 1'b0;
assign COL[19045] = 1'b0;
assign COL[19046] = 1'b0;
assign COL[19047] = 1'b0;
assign COL[19048] = 1'b0;
assign COL[19049] = 1'b0;
assign COL[19050] = 1'b0;
assign COL[19051] = 1'b0;
assign COL[19052] = 1'b0;
assign COL[19053] = 1'b0;
assign COL[19054] = 1'b0;
assign COL[19055] = 1'b0;
assign COL[19056] = 1'b0;
assign COL[19057] = 1'b0;
assign COL[19058] = 1'b0;
assign COL[19059] = 1'b0;
assign COL[19060] = 1'b0;
assign COL[19061] = 1'b0;
assign COL[19062] = 1'b0;
assign COL[19063] = 1'b0;
assign COL[19064] = 1'b0;
assign COL[19065] = 1'b0;
assign COL[19066] = 1'b0;
assign COL[19067] = 1'b0;
assign COL[19068] = 1'b0;
assign COL[19069] = 1'b0;
assign COL[19070] = 1'b0;
assign COL[19071] = 1'b0;
assign COL[19072] = 1'b0;
assign COL[19073] = 1'b0;
assign COL[19074] = 1'b0;
assign COL[19075] = 1'b0;
assign COL[19076] = 1'b0;
assign COL[19077] = 1'b0;
assign COL[19078] = 1'b0;
assign COL[19079] = 1'b0;
assign COL[19080] = 1'b0;
assign COL[19081] = 1'b0;
assign COL[19082] = 1'b0;
assign COL[19083] = 1'b0;
assign COL[19084] = 1'b0;
assign COL[19085] = 1'b0;
assign COL[19086] = 1'b0;
assign COL[19087] = 1'b0;
assign COL[19088] = 1'b0;
assign COL[19089] = 1'b0;
assign COL[19090] = 1'b0;
assign COL[19091] = 1'b0;
assign COL[19092] = 1'b0;
assign COL[19093] = 1'b0;
assign COL[19094] = 1'b0;
assign COL[19095] = 1'b0;
assign COL[19096] = 1'b0;
assign COL[19097] = 1'b0;
assign COL[19098] = 1'b0;
assign COL[19099] = 1'b0;
assign COL[19100] = 1'b0;
assign COL[19101] = 1'b0;
assign COL[19102] = 1'b0;
assign COL[19103] = 1'b0;
assign COL[19104] = 1'b0;
assign COL[19105] = 1'b0;
assign COL[19106] = 1'b0;
assign COL[19107] = 1'b0;
assign COL[19108] = 1'b0;
assign COL[19109] = 1'b0;
assign COL[19110] = 1'b0;
assign COL[19111] = 1'b0;
assign COL[19112] = 1'b0;
assign COL[19113] = 1'b0;
assign COL[19114] = 1'b0;
assign COL[19115] = 1'b0;
assign COL[19116] = 1'b0;
assign COL[19117] = 1'b0;
assign COL[19118] = 1'b0;
assign COL[19119] = 1'b0;
assign COL[19120] = 1'b0;
assign COL[19121] = 1'b0;
assign COL[19122] = 1'b0;
assign COL[19123] = 1'b0;
assign COL[19124] = 1'b0;
assign COL[19125] = 1'b0;
assign COL[19126] = 1'b0;
assign COL[19127] = 1'b0;
assign COL[19128] = 1'b0;
assign COL[19129] = 1'b0;
assign COL[19130] = 1'b0;
assign COL[19131] = 1'b0;
assign COL[19132] = 1'b0;
assign COL[19133] = 1'b0;
assign COL[19134] = 1'b0;
assign COL[19135] = 1'b0;
assign COL[19136] = 1'b0;
assign COL[19137] = 1'b0;
assign COL[19138] = 1'b0;
assign COL[19139] = 1'b0;
assign COL[19140] = 1'b0;
assign COL[19141] = 1'b0;
assign COL[19142] = 1'b0;
assign COL[19143] = 1'b0;
assign COL[19144] = 1'b0;
assign COL[19145] = 1'b0;
assign COL[19146] = 1'b0;
assign COL[19147] = 1'b0;
assign COL[19148] = 1'b0;
assign COL[19149] = 1'b0;
assign COL[19150] = 1'b0;
assign COL[19151] = 1'b0;
assign COL[19152] = 1'b0;
assign COL[19153] = 1'b0;
assign COL[19154] = 1'b0;
assign COL[19155] = 1'b0;
assign COL[19156] = 1'b0;
assign COL[19157] = 1'b0;
assign COL[19158] = 1'b0;
assign COL[19159] = 1'b0;
assign COL[19160] = 1'b0;
assign COL[19161] = 1'b0;
assign COL[19162] = 1'b0;
assign COL[19163] = 1'b0;
assign COL[19164] = 1'b0;
assign COL[19165] = 1'b0;
assign COL[19166] = 1'b0;
assign COL[19167] = 1'b0;
assign COL[19168] = 1'b0;
assign COL[19169] = 1'b0;
assign COL[19170] = 1'b0;
assign COL[19171] = 1'b0;
assign COL[19172] = 1'b0;
assign COL[19173] = 1'b0;
assign COL[19174] = 1'b0;
assign COL[19175] = 1'b0;
assign COL[19176] = 1'b0;
assign COL[19177] = 1'b0;
assign COL[19178] = 1'b0;
assign COL[19179] = 1'b0;
assign COL[19180] = 1'b0;
assign COL[19181] = 1'b0;
assign COL[19182] = 1'b0;
assign COL[19183] = 1'b0;
assign COL[19184] = 1'b0;
assign COL[19185] = 1'b0;
assign COL[19186] = 1'b0;
assign COL[19187] = 1'b0;
assign COL[19188] = 1'b0;
assign COL[19189] = 1'b0;
assign COL[19190] = 1'b0;
assign COL[19191] = 1'b0;
assign COL[19192] = 1'b0;
assign COL[19193] = 1'b0;
assign COL[19194] = 1'b0;
assign COL[19195] = 1'b0;
assign COL[19196] = 1'b0;
assign COL[19197] = 1'b0;
assign COL[19198] = 1'b0;
assign COL[19199] = 1'b0;
assign COL[19200] = 1'b0;


	
	assign location = (x + 1 + (160 * y));	
	assign out = (x > 7'b1001101 && x < 7'b1011001 && y > 7'b0000110 && y < 7'b0010000) ? 2'b10: COL[location];
	


 
endmodule